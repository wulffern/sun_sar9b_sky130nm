magic
tech sky130B
magscale 1 2
timestamp 1708642800
<< checkpaint >>
rect 0 0 2520 704
<< locali >>
rect 864 54 1032 122
rect 1032 54 1656 122
rect 1032 54 1100 122
rect 864 582 1032 650
rect 1032 582 1656 650
rect 1032 582 1100 650
rect 864 406 1032 474
rect 1032 406 1656 474
rect 1032 406 1100 474
rect 398 142 466 386
rect 432 494 600 562
rect 600 54 864 122
rect 600 54 668 562
rect 2088 142 2256 210
rect 2088 494 2256 562
rect 2256 142 2324 562
rect 830 230 898 298
rect 830 406 898 474
rect 1622 230 1690 298
rect 1622 406 1690 474
rect 1980 142 2196 210
rect 1548 406 1764 474
rect 756 582 972 650
<< poly >>
rect 324 158 2196 194
<< m3 >>
rect 1656 230 1824 298
rect 1824 318 2088 386
rect 1824 230 1892 386
rect 1548 0 1732 704
rect 756 0 940 704
rect 1548 0 1732 704
rect 756 0 940 704
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 176
box 0 176 1260 528
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_PCHDL MP0 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1_DMY 
transform 1 0 1260 0 1 176
box 1260 176 2520 528
use SUNSAR_PCHDL MP2 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 230
box 1548 230 1732 298
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 1980 0 1 318
box 1980 318 2164 386
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 1548 0 1 230
box 1548 230 1732 298
use SUNSAR_cut_M1M4_2x1 xcut3 
transform 1 0 756 0 1 230
box 756 230 940 298
use SUNSAR_cut_M1M4_2x1 xcut4 
transform 1 0 756 0 1 230
box 756 230 940 298
<< labels >>
flabel locali s 1980 142 2196 210 0 FreeSans 400 0 0 0 C
port 1 nsew signal bidirectional
flabel locali s 1548 406 1764 474 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 756 582 972 650 0 FreeSans 400 0 0 0 A
port 2 nsew signal bidirectional
flabel m3 s 1548 0 1732 704 0 FreeSans 400 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel m3 s 756 0 940 704 0 FreeSans 400 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 704
<< end >>
