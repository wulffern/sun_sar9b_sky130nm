magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 1260 704
<< locali >>
rect 811 291 845 413
rect 811 467 845 589
rect 432 115 516 149
rect 432 291 516 325
rect 432 379 516 413
rect 516 115 550 413
rect 710 203 828 237
rect 432 643 710 677
rect 710 203 744 677
rect 828 27 912 61
rect 912 599 1044 633
rect 912 27 946 633
rect 378 27 882 61
rect 1206 66 1314 110
rect -54 66 54 110
rect 162 423 270 457
rect 162 247 270 281
rect 990 71 1098 105
rect 162 71 270 105
rect 774 203 882 237
<< poly >>
rect 162 255 1098 273
rect 162 431 1098 449
rect 162 607 1098 625
<< m3 >>
rect 774 0 874 704
rect 378 0 478 704
rect 774 0 874 704
rect 378 0 478 704
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 176
box 0 176 630 352
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 352
box 0 352 630 528
use SUNSAR_NCHDL MN3 
transform 1 0 0 0 1 528
box 0 528 630 704
use SUNSAR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNSAR_PCHDL MP1 
transform 1 0 630 0 1 176
box 630 176 1260 352
use SUNSAR_PCHDL MP2 
transform 1 0 630 0 1 352
box 630 352 1260 528
use SUNSAR_PCHDL MP3 
transform 1 0 630 0 1 528
box 630 528 1260 704
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 115
box 774 115 874 153
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 643
box 774 643 874 681
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 203
box 378 203 478 241
use SUNSAR_cut_M1M4_2x1 xcut3 
transform 1 0 378 0 1 467
box 378 467 478 505
use SUNSAR_cut_M1M4_2x1 xcut4 
transform 1 0 378 0 1 555
box 378 555 478 593
<< labels >>
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel locali s 162 423 270 457 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 990 71 1098 105 0 FreeSans 400 0 0 0 RST_N
port 5 nsew signal bidirectional
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 EN
port 3 nsew signal bidirectional
flabel locali s 774 203 882 237 0 FreeSans 400 0 0 0 ENO
port 4 nsew signal bidirectional
flabel m3 s 774 0 874 704 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 378 0 478 704 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 704
<< end >>
