magic
tech sky130A
magscale 1 2
timestamp 1708902000
<< checkpaint >>
rect 0 0 7272 4800
<< m3 >>
rect -20 760 3672 828
rect -20 1720 3672 1788
rect -20 2680 3672 2748
rect -20 3640 3672 3708
rect -20 4600 3672 4668
rect -20 760 48 4668
rect 3672 -40 7296 28
rect 3672 920 7296 988
rect 3672 1880 7296 1948
rect 3672 2840 7296 2908
rect 3672 3800 7296 3868
rect 7296 -40 7364 3868
rect 108 2680 7236 2760
rect 108 -40 7236 40
use SUNSAR_CAP_BSSW_CV XCAPB0 
transform 1 0 0 0 1 0
box 0 0 7272 960
use SUNSAR_CAP_BSSW_CV XCAPB1 
transform 1 0 0 0 1 960
box 0 960 7272 1920
use SUNSAR_CAP_BSSW_CV XCAPB2 
transform 1 0 0 0 1 1920
box 0 1920 7272 2880
use SUNSAR_CAP_BSSW_CV XCAPB3 
transform 1 0 0 0 1 2880
box 0 2880 7272 3840
use SUNSAR_CAP_BSSW_CV XCAPB4 
transform 1 0 0 0 1 3840
box 0 3840 7272 4800
<< labels >>
flabel m3 s 108 2680 7236 2760 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel m3 s 108 -40 7236 40 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 7272 4800
<< end >>
