magic
tech sky130B
magscale 1 2
timestamp 1672527600
<< checkpaint >>
rect 0 0 76 200
<< m1 >>
rect 0 0 68 184
<< v1 >>
rect 6 12 62 68
rect 6 116 62 172
<< m2 >>
rect 0 0 76 200
<< labels >>
<< end >>
