magic
tech sky130A
timestamp 1708968222
<< locali >>
rect 10296 1303 10428 1337
rect 10394 1239 10428 1303
rect 10394 1205 10488 1239
rect 10458 1171 10512 1205
rect 0 -106 11340 -72
rect 0 -250 11340 -158
rect 0 -394 11340 -302
<< metal1 >>
rect 10296 1567 10630 1601
rect 10296 951 10414 985
rect 10380 457 10414 951
rect 10596 501 10630 1567
rect 10512 467 10630 501
rect 10296 423 10414 457
rect 10380 325 10414 423
rect 10380 291 10512 325
rect 199 -106 233 281
rect 2287 -106 2321 281
rect 2719 -106 2753 281
rect 4807 -106 4841 281
rect 5239 -106 5273 281
rect 7327 -106 7361 281
rect 7759 -106 7793 281
rect 9847 -106 9881 281
<< metal2 >>
rect 378 1990 486 2024
rect 2034 1990 2142 2024
rect 2898 1990 3006 2024
rect 4554 1990 4662 2024
rect 5418 1990 5526 2024
rect 7074 1990 7182 2024
rect 7938 1990 8046 2024
rect 9594 1990 9702 2024
rect 10458 1990 10566 2024
rect 415 1875 449 1990
rect 2071 1875 2105 1990
rect 2935 1875 2969 1990
rect 4591 1875 4625 1990
rect 5455 1875 5489 1990
rect 7111 1875 7145 1990
rect 7975 1875 8009 1990
rect 9631 1875 9665 1990
rect 10495 1963 10529 1990
rect 10512 1787 11340 1821
rect 10178 1479 10296 1513
rect 10178 897 10212 1479
rect 10512 1347 11340 1381
rect 10512 1171 11340 1205
rect 10178 863 10296 897
rect 10178 765 10212 863
rect 10178 731 10512 765
rect 199 -360 233 633
rect 2287 -360 2321 633
rect 2719 -360 2753 633
rect 4807 -360 4841 633
rect 5239 -360 5273 633
rect 7327 -360 7361 633
rect 7759 -360 7793 633
rect 9847 -360 9881 633
rect 162 -394 270 -360
rect 2250 -394 2358 -360
rect 2682 -394 2790 -360
rect 4770 -394 4878 -360
rect 5202 -394 5310 -360
rect 7290 -394 7398 -360
rect 7722 -394 7830 -360
rect 9810 -394 9918 -360
<< metal3 >>
rect 10242 1990 10414 2024
rect 378 -250 470 1936
rect 774 -394 866 1936
rect 1654 -394 1746 1936
rect 2050 -250 2142 1936
rect 2898 -250 2990 1936
rect 3294 -394 3386 1936
rect 4174 -394 4266 1936
rect 4570 -250 4662 1936
rect 5418 -250 5510 1936
rect 5814 -394 5906 1936
rect 6694 -394 6786 1936
rect 7090 -250 7182 1936
rect 7938 -250 8030 1936
rect 8334 -394 8426 1936
rect 9214 -394 9306 1936
rect 9610 -250 9702 1936
rect 10380 633 10414 1990
rect 10296 599 10414 633
rect 10178 247 10296 281
rect 10178 -360 10212 247
rect 10458 -250 10550 176
rect 10178 -394 10350 -360
rect 10854 -394 10946 176
use SUNSAR_IVX1_CV  SUNSAR_IVX1_CV_0
timestamp 1708968222
transform 1 0 10080 0 1 176
box -90 -66 1350 242
use SUNSAR_TAPCELLB_CV  XA1
timestamp 1708968222
transform 1 0 10080 0 1 0
box -90 -66 1350 242
use SUNSAR_TIEL_CV  XA2
timestamp 1708968222
transform 1 0 10080 0 1 1848
box -90 -66 1350 242
use SUNSAR_IVX1_CV  XA3
timestamp 1708968222
transform 1 0 10080 0 1 352
box -90 -66 1350 242
use SUNSAR_BFX1_CV  XA4
timestamp 1708902000
transform 1 0 10080 0 1 528
box -90 -66 1350 330
use SUNSAR_IVX1_CV  XA5a
timestamp 1708968222
transform 1 0 10080 0 1 1232
box -90 -66 1350 242
use SUNSAR_ORX1_CV  XA5
timestamp 1708968222
transform 1 0 10080 0 1 792
box -90 -66 1350 506
use SUNSAR_ANX1_CV  XA6
timestamp 1708968222
transform 1 0 10080 0 1 1408
box -90 -66 1350 506
use SUNSAR_DFQNX1_CV  XB07
timestamp 1708968222
transform 1 0 0 0 1 0
box -90 -66 1350 2002
use SUNSAR_DFQNX1_CV  XC08
timestamp 1708968222
transform -1 0 2520 0 1 0
box -90 -66 1350 2002
use SUNSAR_cut_M1M2_2x1  xcut0
timestamp 1708902000
transform 1 0 170 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut1
timestamp 1708902000
transform 1 0 170 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut2
timestamp 1708902000
transform 1 0 2258 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut3
timestamp 1708902000
transform 1 0 2258 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut4
timestamp 1708902000
transform 1 0 2690 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut5
timestamp 1708902000
transform 1 0 2690 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut6
timestamp 1708902000
transform 1 0 4778 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut7
timestamp 1708902000
transform 1 0 4778 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut8
timestamp 1708902000
transform 1 0 5210 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut9
timestamp 1708902000
transform 1 0 5210 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut10
timestamp 1708902000
transform 1 0 7298 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut11
timestamp 1708902000
transform 1 0 7298 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut12
timestamp 1708902000
transform 1 0 7730 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut13
timestamp 1708902000
transform 1 0 7730 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut14
timestamp 1708902000
transform 1 0 9818 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut15
timestamp 1708902000
transform 1 0 9818 0 1 -106
box 0 0 92 34
use SUNSAR_cut_M1M4_2x2  xcut16
timestamp 1708902000
transform 1 0 378 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut17
timestamp 1708902000
transform 1 0 2050 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut18
timestamp 1708902000
transform 1 0 2898 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut19
timestamp 1708902000
transform 1 0 4570 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut20
timestamp 1708902000
transform 1 0 5418 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut21
timestamp 1708902000
transform 1 0 7090 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut22
timestamp 1708902000
transform 1 0 7938 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut23
timestamp 1708902000
transform 1 0 9610 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut24
timestamp 1708902000
transform 1 0 10458 0 1 -250
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut25
timestamp 1708902000
transform 1 0 774 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut26
timestamp 1708902000
transform 1 0 1654 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut27
timestamp 1708902000
transform 1 0 3294 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut28
timestamp 1708902000
transform 1 0 4174 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut29
timestamp 1708902000
transform 1 0 5814 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut30
timestamp 1708902000
transform 1 0 6694 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut31
timestamp 1708902000
transform 1 0 8334 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut32
timestamp 1708902000
transform 1 0 9214 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M4_2x2  xcut33
timestamp 1708902000
transform 1 0 10854 0 1 -394
box 0 0 92 92
use SUNSAR_cut_M1M2_2x1  xcut34
timestamp 1708902000
transform 1 0 10242 0 1 423
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut35
timestamp 1708902000
transform 1 0 10458 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut36
timestamp 1708902000
transform 1 0 10242 0 1 951
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut37
timestamp 1708902000
transform 1 0 10458 0 1 467
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut38
timestamp 1708902000
transform 1 0 10242 0 1 1567
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut39
timestamp 1708902000
transform 1 0 10258 0 1 863
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut40
timestamp 1708902000
transform 1 0 10474 0 1 731
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut41
timestamp 1708902000
transform 1 0 10258 0 1 1479
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut42
timestamp 1708902000
transform 1 0 170 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut43
timestamp 1708902000
transform 1 0 2258 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut44
timestamp 1708902000
transform 1 0 2690 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut45
timestamp 1708902000
transform 1 0 4778 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut46
timestamp 1708902000
transform 1 0 5210 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut47
timestamp 1708902000
transform 1 0 7298 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut48
timestamp 1708902000
transform 1 0 7730 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut49
timestamp 1708902000
transform 1 0 9818 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut50
timestamp 1708902000
transform 1 0 9602 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut51
timestamp 1708902000
transform 1 0 7946 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut52
timestamp 1708902000
transform 1 0 7082 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut53
timestamp 1708902000
transform 1 0 5426 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut54
timestamp 1708902000
transform 1 0 4562 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut55
timestamp 1708902000
transform 1 0 2906 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut56
timestamp 1708902000
transform 1 0 2042 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut57
timestamp 1708902000
transform 1 0 386 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut58
timestamp 1708902000
transform 1 0 10458 0 1 1171
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut59
timestamp 1708902000
transform 1 0 10458 0 1 1347
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut60
timestamp 1708902000
transform 1 0 10458 0 1 1787
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut61
timestamp 1708902000
transform 1 0 10242 0 1 599
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut62
timestamp 1708902000
transform 1 0 10466 0 1 1963
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut63
timestamp 1708902000
transform 1 0 10258 0 1 247
box 0 0 92 34
use SUNSAR_DFQNX1_CV  XD09
timestamp 1708968222
transform 1 0 2520 0 1 0
box -90 -66 1350 2002
use SUNSAR_DFQNX1_CV  XE10
timestamp 1708968222
transform -1 0 5040 0 1 0
box -90 -66 1350 2002
use SUNSAR_DFQNX1_CV  XF11
timestamp 1708968222
transform 1 0 5040 0 1 0
box -90 -66 1350 2002
use SUNSAR_DFQNX1_CV  XG12
timestamp 1708968222
transform -1 0 7560 0 1 0
box -90 -66 1350 2002
use SUNSAR_DFQNX1_CV  XH13
timestamp 1708968222
transform 1 0 7560 0 1 0
box -90 -66 1350 2002
use SUNSAR_DFQNX1_CV  XI14
timestamp 1708968222
transform -1 0 10080 0 1 0
box -90 -66 1350 2002
<< labels >>
flabel locali s 0 -106 11340 -72 0 FreeSans 200 0 0 0 DONE
port 22 nsew signal bidirectional
flabel locali s 0 -250 11340 -158 0 FreeSans 200 0 0 0 AVSS
port 24 nsew signal bidirectional
flabel locali s 0 -394 11340 -302 0 FreeSans 200 0 0 0 AVDD
port 23 nsew signal bidirectional
flabel metal3 s 10242 1990 10350 2024 0 FreeSans 200 0 0 0 CKS
port 1 nsew signal bidirectional
flabel metal3 s 10242 -394 10350 -360 0 FreeSans 200 0 0 0 ENABLE
port 2 nsew signal bidirectional
flabel metal2 s 11232 1171 11340 1205 0 FreeSans 200 0 0 0 CK_SAMPLE
port 3 nsew signal bidirectional
flabel metal2 s 11232 1787 11340 1821 0 FreeSans 200 0 0 0 CK_SAMPLE_BSSW
port 4 nsew signal bidirectional
flabel metal2 s 11232 1347 11340 1381 0 FreeSans 200 0 0 0 EN
port 5 nsew signal bidirectional
flabel metal2 s 162 -394 270 -360 0 FreeSans 200 0 0 0 D<7>
port 6 nsew signal bidirectional
flabel metal2 s 2250 -394 2358 -360 0 FreeSans 200 0 0 0 D<6>
port 7 nsew signal bidirectional
flabel metal2 s 2682 -394 2790 -360 0 FreeSans 200 0 0 0 D<5>
port 8 nsew signal bidirectional
flabel metal2 s 4770 -394 4878 -360 0 FreeSans 200 0 0 0 D<4>
port 9 nsew signal bidirectional
flabel metal2 s 5202 -394 5310 -360 0 FreeSans 200 0 0 0 D<3>
port 10 nsew signal bidirectional
flabel metal2 s 7290 -394 7398 -360 0 FreeSans 200 0 0 0 D<2>
port 11 nsew signal bidirectional
flabel metal2 s 7722 -394 7830 -360 0 FreeSans 200 0 0 0 D<1>
port 12 nsew signal bidirectional
flabel metal2 s 9810 -394 9918 -360 0 FreeSans 200 0 0 0 D<0>
port 13 nsew signal bidirectional
flabel metal2 s 378 1990 486 2024 0 FreeSans 200 0 0 0 DO<7>
port 14 nsew signal bidirectional
flabel metal2 s 2034 1990 2142 2024 0 FreeSans 200 0 0 0 DO<6>
port 15 nsew signal bidirectional
flabel metal2 s 2898 1990 3006 2024 0 FreeSans 200 0 0 0 DO<5>
port 16 nsew signal bidirectional
flabel metal2 s 4554 1990 4662 2024 0 FreeSans 200 0 0 0 DO<4>
port 17 nsew signal bidirectional
flabel metal2 s 5418 1990 5526 2024 0 FreeSans 200 0 0 0 DO<3>
port 18 nsew signal bidirectional
flabel metal2 s 7074 1990 7182 2024 0 FreeSans 200 0 0 0 DO<2>
port 19 nsew signal bidirectional
flabel metal2 s 7938 1990 8046 2024 0 FreeSans 200 0 0 0 DO<1>
port 20 nsew signal bidirectional
flabel metal2 s 9594 1990 9702 2024 0 FreeSans 200 0 0 0 DO<0>
port 21 nsew signal bidirectional
flabel metal2 s 10458 1990 10566 2024 0 FreeSans 200 0 0 0 TIE_L
port 25 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 -394 11340 2024
<< end >>
