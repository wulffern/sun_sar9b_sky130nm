magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect 0 0 8712 5280
<< m3 >>
rect -40 836 4392 912
rect -40 1892 4392 1968
rect -40 2948 4392 3024
rect -40 4004 4392 4080
rect -40 5060 4392 5136
rect -40 836 36 5136
rect 4392 -44 8748 32
rect 4392 1012 8748 1088
rect 4392 2068 8748 2144
rect 4392 3124 8748 3200
rect 4392 4180 8748 4256
rect 8748 -44 8824 4256
rect 108 2948 8676 3036
rect 108 -44 8676 44
use SUNSAR_CAP_BSSW_CV XCAPB0 
transform 1 0 0 0 1 0
box 0 0 8712 1056
use SUNSAR_CAP_BSSW_CV XCAPB1 
transform 1 0 0 0 1 1056
box 0 1056 8712 2112
use SUNSAR_CAP_BSSW_CV XCAPB2 
transform 1 0 0 0 1 2112
box 0 2112 8712 3168
use SUNSAR_CAP_BSSW_CV XCAPB3 
transform 1 0 0 0 1 3168
box 0 3168 8712 4224
use SUNSAR_CAP_BSSW_CV XCAPB4 
transform 1 0 0 0 1 4224
box 0 4224 8712 5280
<< labels >>
flabel m3 s 108 2948 8676 3036 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel m3 s 108 -44 8676 44 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 8712 0 5280
<< end >>
