* NGSPICE file created from SUNSAR_SAR9B_CV.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW
+ VREF AVDD AVSS
*.subckt SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4>
*+ D<3> D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
X0 XA20.XA10.A CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 XA20.XA11.MP1.S CK_SAMPLE AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 VREF XA4.XA1.CHL_OP XA4.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X3 XA6.XA6.MP3.S D<2> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X4 SAR_IN XB2.CKN XB2.XA3.B AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X5 XA7.XA10.A XA7.XA6.Y XA7.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R0 XDAC1.XC128a<1>.XRES2.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R1 XDAC1.XC1.XRES4.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X6 AVDD XA7.XA6.Y XA7.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X7 XA20.XA4.MP0.S SARN XA20.XA4.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X8 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=134.8596 ps=707.66 w=1.08 l=0.18
X9 XA6.CP0 XA6.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R2 XDAC1.XC64a<0>.XRES1A.B XA1.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X10 XA2.XA1.XA5.MP2.S EN XA2.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X11 XA0.CMP_ON XA20.XA2.CO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 XDAC1.XC32a<0>.XRES1B.B D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X12 SAR_IN XB2.XA3.MP0.S XB2.XA3.B AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X13 XA6.XA10.Y XA6.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X14 XA0.CMP_ON XA20.XA2.CO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X15 XA6.XA2.A EN XA6.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X16 XA2.XA11.Y XA2.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X17 AVSS XA5.CEO XA6.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 XA6.XA6.MP1.S XA6.CN0 XA6.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X19 XA20.XA2.N2 SARP XA20.XA2.N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X20 D<0> XA8.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 XA6.XA1.XA1.MP3.S XA0.CMP_OP XA6.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 XA20.XA2.CO XA20.XA1.CK AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X23 XA2.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R4 XDAC1.X16ab.XRES2.B D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R5 XDAC1.XC64b<1>.XRES2.B D<7> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X24 XA6.XA6.Y CK_SAMPLE XA6.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X25 VREF XA6.CN1 D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X26 XA2.CP0 XA2.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 XA1.XA9.MN1.S XA1.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R6 XA0.CN0 XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X28 XA1.XA10.A XA1.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X29 XA20.XA4.MP0.S SARN XA20.XA4.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X30 XA0.CMP_ON XA20.XA2.CO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X31 XA0.CMP_ON XA20.XA2.CO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X32 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X33 AVSS XA6.XA1.CHL_OP XA6.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X34 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=203.8716 ps=1.06874k w=1.08 l=0.18
X35 XA6.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X36 XA2.XA10.Y XA2.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 XA2.XA2.A XA1.ENO XA2.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X38 XA1.CN0 XA1.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R7 XA1.CN0 XDAC2.XC64a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X39 XA20.XA2.N2 SARP XA20.XA2.N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X40 XA1.CN0 XA1.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X41 XA20.XA2.N2 XA20.XA1.CK AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X42 XA2.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 AVSS XA5.CP0 XA5.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 VREF XA5.CP0 XA5.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 AVSS XA0.CMP_OP XA2.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X46 D<7> XA1.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X47 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X48 AVSS CK_SAMPLE XA6.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X49 D<7> XA1.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X50 AVSS XA2.CN1 D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X51 AVSS XA5.CN1 D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R8 m3_830_1080# XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X52 VREF XA5.CN1 D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X53 AVSS XA3.XA2.A XA3.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R9 XDAC1.XC32a<0>.XRES2.B D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X54 XA20.XA1.MP0.S SARP XA20.XA1.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X55 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X56 XA1.XA1.XA4.MN2.S XA1.XA1.XA4.LCK_N XA1.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X57 AVSS XA0.XA2.A D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X58 VREF XA3.XA2.A XA3.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X59 XA1.XA1.XA4.MP2.S EN XA1.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X60 XA0.CP1 D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X61 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X62 XA2.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X63 XA8.XA1.XA5.MP2.S EN XA8.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X64 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X65 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X66 XA8.XA11.Y XA8.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X67 AVSS XA5.CP0 XA5.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X68 XA3.DONE XA3.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 VREF XA5.CP0 XA5.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X70 AVSS XA1.XA2.A XA1.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X71 XA3.DONE XA3.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X72 VREF XA1.XA2.A XA1.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X73 XA0.DONE XA0.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R10 m3_16526_2200# XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X74 XA8.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X75 XA20.XA1.MP0.S XA20.XA1.CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X76 XA3.CN0 XA3.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X77 AVDD XA20.XA1.CKN XA20.XA1.MP0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X78 XA4.XA11.MP1.S XA4.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X79 XA0.CN0 XA0.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 XA3.CN0 XA3.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 XA4.CEIN XA3.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 XA8.CP0 XA8.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 AVSS XA7.XA2.A XA7.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R11 XDAC1.XC0.XRES8.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X84 XA4.CEIN XA3.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 VREF XA7.XA2.A XA7.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X86 XA0.CEO XA0.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X87 XA4.XA6.MP3.S D<4> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X88 XA8.XA10.Y XA8.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X89 XA5.XA10.A XA5.XA6.Y XA5.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X90 XA1.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X91 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X92 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X93 AVDD XA5.XA6.Y XA5.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X94 XA3.XA8.A XA4.EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X95 XA1.XA1.XA1.MP2.S XA0.CMP_ON XA1.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X96 XA8.XA2.A XA7.ENO XA8.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X97 XA0.XA8.A XA0.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X98 XA3.XA8.A XA4.EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X99 XA4.CP0 XA4.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X100 XA7.DONE XA7.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X101 XA8.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 XA0.XA1.XA5.MP2.S EN XA0.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X103 SAR_IP XB1.CKN XB1.XA3.B AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X104 AVSS XA0.CMP_OP XA8.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 XA7.DONE XA7.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X106 AVSS XA3.XA1.CHL_OP XA3.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X107 XA4.XA10.Y XA4.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X108 AVSS XA0.XA1.CHL_OP XA0.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X109 VREF XA3.XA1.CHL_OP XA3.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X110 XA4.XA2.A EN XA4.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X111 AVSS XA8.CN1 D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R12 XDAC1.XC64a<0>.XRES2.B XA1.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X112 XA7.CN0 XA7.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 XA2.XA1.CHL_OP EN XA2.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X114 AVSS XA4.CEIN XA4.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X115 XA4.XA6.MP1.S XA4.CN0 XA4.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X116 XA7.CN0 XA7.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 XA6.XA10.A XA6.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R13 XA0.CN0 XDAC2.XC128b<2>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X118 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X119 XA4.XA1.XA1.MP3.S XA0.CMP_OP XA4.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X120 XA7.CEO XA7.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X121 XA1.XA1.XA1.MN2.S XA0.ENO XA1.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X122 XA8.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X123 XA7.CEO XA7.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X124 XA20.XA1.CK XA20.XA1.CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X125 SAR_IP XB1.M1.G SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X126 AVDD EN XA1.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X127 XA20.XA1.CK XA20.XA1.CKN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X128 XA4.XA6.Y CK_SAMPLE XA4.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X129 VREF XA4.CN1 D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X130 XA6.CN0 XA6.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X131 XA7.XA8.A XA7.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R14 XDAC1.X16ab.XRES4.B D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R15 XDAC1.XC64b<1>.XRES4.B D<7> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X132 XA7.XA8.A XA7.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X133 XA20.XA2.N1 SARN XA20.XA3.N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X134 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X135 AVSS XA4.XA1.CHL_OP XA4.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X136 AVDD XA20.XA2.CO XA20.XA2.VMR AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X137 XA4.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X138 D<2> XA6.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X139 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X140 AVSS XA7.XA1.CHL_OP XA7.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R16 XDAC1.XC0.XRES1A.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X141 XA2.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X142 VREF XA7.XA1.CHL_OP XA7.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 XA0.CMP_OP XA20.XA2.VMR AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X144 XA0.CMP_OP XA20.XA2.VMR AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X145 XB2.XA1.Y XB2.XA1.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X146 XA6.XA1.XA4.MP2.S EN XA6.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X147 XA2.XA9.MN1.S XA2.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X148 SAR_IN XB1.TIE_L SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X149 AVSS CK_SAMPLE XA4.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X150 AVDD XA20.XA1.CK XA20.XA1.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X151 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X152 XA2.CN0 XA2.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X153 XB2.XA1.MP0.G XB2.XA1.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X154 AVSS XA6.CP0 XA6.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X155 VREF XA6.XA2.A XA6.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X156 D<6> XA2.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X158 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X159 XA20.XA2.VMR XA20.XA2.CO XA20.XA3.N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R17 XB2.XA4.GNG m3_23222_3960# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X160 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X161 AVDD XA20.XA2.CO XA20.XA2.VMR AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X162 AVSS XA6.CN1 D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R18 XDAC1.XC128b<2>.XRES1A.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R19 XB1.XA3.B m3_7598_4120# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X163 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X164 SAR_IN XB1.TIE_L SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X165 XA8.XA1.CHL_OP EN XA8.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X166 XA2.XA1.XA4.MN2.S XA2.XA1.XA4.LCK_N XA2.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X167 XA1.CP0 XA1.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X168 XA1.CP0 XA1.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X169 XA1.CN1 XA1.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X170 XA6.XA1.XA1.MP2.S XA0.CMP_ON XA6.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 AVSS XA6.CP0 XA6.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X172 XA1.CN1 XA1.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 XA20.XA2.N1 XA20.XA1.CK AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X174 AVDD XA20.XA1.CK XA20.XA2.N1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X175 AVSS XA2.XA2.A XA2.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X176 AVSS XA5.XA2.A XA5.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X177 SAR_IP XB1.M1.G SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X178 VREF XA5.XA2.A XA5.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X179 XA1.ENO XA1.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 AVDD XA1.XA1.XA1.MP3.G XA1.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X181 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X182 XA3.XA11.Y XA3.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X183 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X185 XA8.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X186 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X187 XA3.XA11.MP1.S XA3.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X188 XA0.XA11.Y XA0.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X189 XA8.XA9.MN1.S XA8.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 XA5.DONE XA5.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X191 XA5.DONE XA5.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 XA3.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X193 XA3.XA6.MP3.S D<5> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X194 AVDD EN XA6.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X195 XA6.XA10.A XA6.XA6.Y XA6.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X196 XA0.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X197 XA2.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X198 XA5.CN0 XA5.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X199 XA8.CN0 XA8.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R20 m3_16526_280# XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X200 XA0.XA1.CHL_OP EN XA0.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X201 XA5.CN0 XA5.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X202 XA3.CP0 XA3.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X203 XA1.CN1 XA1.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 XA4.XA10.A XA4.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X205 XA3.CP0 XA3.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X206 XA1.CN1 XA1.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X207 XA5.CEO XA5.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X208 XA0.CP0 XA0.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R21 D<8> XDAC2.XC128a<1>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R22 XA5.CN0 XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X209 XA5.CEO XA5.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X210 XA3.XA10.Y XA3.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X211 D<0> XA8.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X212 XA3.XA10.Y XA3.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X213 XA3.XA2.A XA2.ENO XA3.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X214 XA1.XA1.XA4.LCK_N XA1.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X215 XA0.XA10.Y XA0.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X216 XA4.CN0 XA4.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X217 XA0.XA2.A EN XA0.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X218 XA3.XA2.A EN XA3.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R23 XA3.CN1 XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X219 XA1.XA1.XA4.LCK_N XA1.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X220 XA5.XA8.A XA5.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X221 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X222 XA7.XA11.Y XA7.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X223 XA5.XA8.A XA5.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X224 XA3.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X225 XA8.XA1.XA4.MN2.S XA8.XA1.XA4.LCK_N XA8.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X226 XA7.XA11.MP1.S XA7.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X227 XA0.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X228 XA3.XA6.MP1.S XA3.CN0 XA3.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R24 XA1.CN1 XDAC2.XC64b<1>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X229 AVSS XA0.CMP_OP XA3.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X230 D<4> XA4.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X231 XA2.XA1.XA1.MN2.S XA1.ENO XA2.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X232 XA3.XA1.XA1.MP3.S XA0.CMP_OP XA3.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X233 AVSS XA0.CMP_OP XA0.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X234 XA7.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X235 AVSS XA5.XA1.CHL_OP XA5.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X236 SAR_IN XB2.M1.G SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X237 XA0.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X238 XA7.XA6.MP3.S D<1> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X239 VREF XA5.XA1.CHL_OP XA5.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X240 AVSS XA3.CN1 D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X241 AVSS D<8> XA0.CP1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X242 VREF XA3.CN1 D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X243 XA4.XA1.XA4.MP2.S EN XA4.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X244 AVSS XA8.XA2.A XA8.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 XA7.CP0 XA7.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X246 XA7.CP0 XA7.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X247 XA3.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X248 XA0.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 XA3.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R25 XA0.CN0 XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R26 D<8> XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X250 XB2.XA4.GNG XB2.CKN XB2.M1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X251 XA7.XA10.Y XA7.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X252 XB1.XA1.Y XB1.XA1.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X253 XA7.XA10.Y XA7.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X254 XA7.XA2.A XA6.ENO XA7.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X255 AVSS XA4.CP0 XA4.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X256 VREF XA4.XA2.A XA4.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X257 XA7.XA2.A EN XA7.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X258 XA6.CP0 XA6.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X259 XA7.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X260 XA7.XA6.MP1.S XA7.CN0 XA7.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R27 D<8> XDAC2.XC128a<1>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R28 XA2.CN1 XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X261 XB2.XA4.MN1.S XB2.CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 AVSS XA0.CMP_OP XA7.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X263 AVSS XA4.CN1 D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X264 XA8.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X265 XA7.XA1.XA1.MP3.S XA0.CMP_OP XA7.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X266 XA6.CN1 XA6.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X267 AVSS XA7.CN1 D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X268 VREF XA7.CN1 D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X269 XA20.XA2.N2 SARP XA20.XA2.N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X270 AVDD XA6.XA1.XA1.MP3.G XA6.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 XA20.XA2.CO XA20.XA2.VMR AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X272 XA4.XA1.XA1.MP2.S XA0.CMP_ON XA4.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X273 XA7.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X274 AVSS XA4.CP0 XA4.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R29 XA0.CN0 XDAC2.XC128b<2>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X275 XA7.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X276 XA2.CP0 XA2.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R30 XA2.CN0 XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X277 XA8.XA1.XA1.MN2.S XA7.ENO XA8.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X278 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X279 XA2.CN1 XA2.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R31 D<8> XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X280 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X281 XA20.XA3.N2 SARN XA20.XA2.N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X282 XA20.XA3.N2 XA20.XA1.CK AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X283 XA6.CN1 XA6.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X284 AVSS XA6.XA2.A XA6.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X285 XA2.XA11.Y XA1.CEO XA2.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X286 XA2.ENO XA2.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 D<7> XA1.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X288 XB1.CKN CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 AVDD EN XA4.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X291 XA4.XA10.A XA4.XA6.Y XA4.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X292 D<7> XA1.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X293 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X294 XA6.XA1.XA4.LCK_N XA6.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X295 XA2.XA6.Y D<6> XA2.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X296 XA6.DONE XA6.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X297 XA20.XA1.MP0.S SARP XA20.XA1.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X298 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X299 VREF XA2.XA1.CHL_OP XA2.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X300 XA6.CN0 XA6.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X301 XA5.XA11.Y XA5.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X302 XA3.XA9.MN1.S XA3.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 XA2.CN1 XA2.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X304 XA5.XA11.MP1.S XA5.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X305 XA3.XA10.A XA3.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X306 XA6.CEO XA6.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X307 XA0.XA9.MN1.S XA0.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X308 XA5.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X309 AVDD XA2.CN0 XA2.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X310 XA5.XA6.MP3.S D<3> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X311 XA3.CN0 XA3.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X312 XA2.XA1.XA4.LCK_N XA2.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X313 XA3.CN0 XA3.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R32 XA1.CN1 XDAC2.XC64b<1>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X314 XA6.XA8.A XA6.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X315 XA0.CN0 XA0.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X316 XA5.CP0 XA5.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X317 XA8.CP0 XA8.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X318 XA5.CP0 XA5.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X319 D<5> XA3.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X320 D<5> XA3.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X321 XA1.XA1.XA5.MP2.S EN XA1.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X322 XA1.XA1.XA5.MN2.S XA1.XA1.XA4.LCK_N XA1.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X323 XA5.XA10.Y XA5.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X324 AVSS XA6.XA1.CHL_OP XA6.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X325 XA0.CP1 D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 XA5.XA10.Y XA5.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X327 XA8.CN1 XA8.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X328 XA5.XA2.A XA4.ENO XA5.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X329 XA5.XA2.A EN XA5.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X330 SAR_IP XB1.TIE_L SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X331 XA3.XA1.XA4.MN2.S XA3.XA1.XA4.LCK_N XA3.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X332 XA4.CP0 XA4.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X333 XA3.XA1.XA4.MP2.S EN XA3.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X334 XA0.XA1.XA4.MN2.S XA0.XA1.XA4.LCK_N XA0.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X335 XA8.XA11.Y XA7.CEO XA8.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X336 XA5.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X337 XB1.XA4.GNG XB1.CKN XB1.M1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X338 XA7.XA9.MN1.S XA7.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X339 XA5.XA6.MP1.S XA5.CN0 XA5.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X340 AVSS XA0.CMP_OP XA5.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X341 XA8.ENO XA8.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X342 XA7.XA10.A XA7.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X343 XA5.XA1.XA1.MP3.S XA0.CMP_OP XA5.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X344 XA4.CN1 XA4.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R33 XB2.XA4.GNG m3_23222_3000# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X345 XA8.XA6.Y D<0> XA8.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X346 XA7.CN0 XA7.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X347 AVSS XA5.CN1 D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X348 XA7.CN0 XA7.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X349 VREF XA5.CN1 D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X350 AVSS XA3.XA2.A XA3.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R34 XA4.CN0 XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X351 AVSS XA0.XA2.A D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X352 VREF XA3.XA2.A XA3.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X353 XB2.XA2.MP0.G XB2.XA2.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X354 AVDD XA4.XA1.XA1.MP3.G XA4.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X355 VREF XA8.XA1.CHL_OP XA8.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X356 D<1> XA7.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SAR_IP XB1.TIE_L SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 XB1.M1.G XB1.XA1.Y XB1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X359 XA5.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X360 D<1> XA7.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X361 XA5.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 XA8.CN1 XA8.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X363 XB1.TIE_L XB2.XA2.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X364 XA7.XA1.XA4.MN2.S XA7.XA1.XA4.LCK_N XA7.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X365 XA7.XA1.XA4.MP2.S EN XA7.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X366 D<2> XA6.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R35 XDAC1.XC1.XRES16.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X367 AVDD XA8.CN0 XA8.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X368 XA3.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X369 XA8.XA1.XA4.LCK_N XA8.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R36 XA3.CN0 XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X370 XA3.XA1.XA1.MP2.S XA0.CMP_ON XA4.EN AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X371 XA0.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X372 AVSS XA4.XA2.A XA4.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X373 XA0.XA11.Y XB1.TIE_L XA0.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X374 XA4.CN1 XA4.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X375 AVSS XA7.XA2.A XA7.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X376 VREF XA7.XA2.A XA7.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X377 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X378 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X379 XA4.XA1.XA4.LCK_N XA4.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X380 XA0.XA6.Y XA0.CP1 XA0.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R37 XDAC1.XC128b<2>.XRES8.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X381 XA4.DONE XA4.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X382 XA20.XA2.N1 SARP XA20.XA2.N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X383 XB2.XA3.B AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X384 AVDD XA20.XA2.VMR XA20.XA2.CO AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X385 VREF XA0.XA1.CHL_OP XA0.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X386 D<6> XA2.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X387 XA3.XA1.XA1.MN2.S XA2.ENO XA3.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X388 AVDD EN XA3.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X389 XA0.XA1.XA1.MN2.S EN XA0.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X390 XA4.CN0 XA4.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R38 XA0.CN0 XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X391 XA7.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X392 XA7.XA1.XA1.MP2.S XA0.CMP_ON XA7.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X393 XA4.CEO XA4.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X394 AVSS XA20.XA2.CO XA0.CMP_ON AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R39 XA1.CN0 XDAC2.XC64a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X395 XB2.XA3.B XB2.CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X396 AVDD XA20.XA2.CO XA0.CMP_ON AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R40 XB1.XA3.B m3_7598_2200# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X397 AVDD XA0.CN0 XA0.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X398 XA6.XA1.XA5.MP2.S EN XA6.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X399 XA4.XA8.A XA4.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X400 XA20.XA2.N1 SARP XA20.XA2.N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X401 XA6.XA11.Y XA6.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X402 AVDD AVDD XA20.XA2.N2 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X403 VREF XA2.CP0 XA2.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R41 XA3.CN1 XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X404 XA6.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X405 AVSS XA4.XA1.CHL_OP XA4.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X406 XA7.XA1.XA1.MN2.S XA6.ENO XA7.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X407 VREF XA2.CN1 D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X408 AVDD EN XA7.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X409 XA1.XA1.CHL_OP XA0.ENO XA1.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X410 XA6.CP0 XA6.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X411 XA1.XA1.CHL_OP EN XA1.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X412 XA5.XA9.MN1.S XA5.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X413 XA2.XA1.XA5.MN2.S XA2.XA1.XA4.LCK_N XA2.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X414 XA5.XA10.A XA5.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 XA6.XA10.Y XA6.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X416 XA6.XA2.A XA5.ENO XA6.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X417 VREF XA2.CP0 XA2.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X418 XA5.CN0 XA5.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X419 XA5.CN0 XA5.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X420 XA3.CP0 XA3.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X421 XA3.CP0 XA3.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X422 XA6.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X423 XA0.CP0 XA0.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X424 D<3> XA5.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X425 D<0> XA8.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X426 AVSS XA0.CMP_OP XA6.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X427 D<3> XA5.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X428 XA3.CN1 XA3.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X429 XA3.CN1 XA3.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X430 XA1.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X431 AVSS XA6.CN1 D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X432 D<8> XA0.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X433 XB1.XA2.MP0.G XB1.XA2.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X434 XA1.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R42 XA0.CN0 XDAC2.XC128b<2>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X435 XA5.XA1.XA4.MN2.S XA5.XA1.XA4.LCK_N XA5.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X436 XA4.EN XA3.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X437 XA5.XA1.XA4.MP2.S EN XA5.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X438 D<4> XA4.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X439 AVDD XA3.XA1.XA1.MP3.G XA3.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X440 XA0.ENO XA0.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X441 XA6.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X442 AVDD XA2.XA6.Y XA2.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X443 XB1.CKN CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R43 m3_16526_3160# XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X444 VREF XA8.CP0 XA8.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X445 XA7.CP0 XA7.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X446 AVSS XA5.XA2.A XA5.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X447 XA20.XA10.MN1.S XA20.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X448 XA7.CP0 XA7.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X449 VREF XA5.XA2.A XA5.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X450 XA20.XA1.CKN XA20.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X451 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X452 VREF XA8.CN1 D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X453 XA7.CN1 XA7.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R44 XDAC1.XC128a<1>.XRES4.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R45 XDAC1.XC32a<0>.XRES4.B D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X454 XA3.CN1 XA3.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X455 XA7.CN1 XA7.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X456 D<8> XA0.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X457 XA3.CN1 XA3.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R46 XDAC1.X16ab.XRES1B.B D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X458 XA7.ENO XA7.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X459 XA8.XA1.XA5.MN2.S XA8.XA1.XA4.LCK_N XA8.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X460 AVDD XA7.XA1.XA1.MP3.G XA7.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X461 XA3.XA1.XA4.LCK_N XA4.EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R47 XDAC1.XC64b<1>.XRES16.B D<7> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X462 XA5.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X463 XA3.XA1.XA4.LCK_N XA4.EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X464 XA0.XA1.XA4.LCK_N XA0.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X465 VREF XA8.CP0 XA8.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X466 XB1.XA3.B AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X467 XA5.XA1.XA1.MP2.S XA0.CMP_ON XA5.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X468 XA4.XA1.XA5.MP2.S EN XA4.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R48 XA0.CN0 XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R49 m3_830_2040# XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X469 XA4.XA11.Y XA4.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R50 XA1.CN0 XDAC2.XC64a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X470 VREF XA0.CP0 XA0.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R51 XDAC1.XC0.XRES1B.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X471 XA6.XA1.CHL_OP EN XA6.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X472 XA7.CN1 XA7.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X473 SAR_IP XB1.XA3.MP0.S XB1.XA3.B AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X474 XA4.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X475 XA7.CN1 XA7.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X476 XA5.XA1.XA1.MN2.S XA4.ENO XA5.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X477 AVDD XA8.XA6.Y XA8.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X478 VREF D<8> XA0.CP1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X479 AVDD EN XA5.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X480 XA7.XA1.XA4.LCK_N XA7.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X481 XA4.CP0 XA4.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R52 XDAC1.XC128a<1>.XRES16.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R53 XDAC1.XC32a<0>.XRES16.B D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R54 XDAC1.XC1.XRES8.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X482 XA7.XA1.XA4.LCK_N XA7.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SAR_IN XB2.M1.G SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X484 AVDD XB1.CKN XB1.XA3.MP0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X485 XA4.XA10.Y XA4.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X486 AVSS XA20.XA2.VMR XA0.CMP_OP AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X487 AVDD XA20.XA2.VMR XA0.CMP_OP AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X488 XA4.XA2.A XA4.EN XA4.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X489 VREF XA0.CP0 XA0.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X490 XA6.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X491 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X492 XA2.XA1.CHL_OP XA1.ENO XA2.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X493 XA4.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R55 XB2.XA4.GNG m3_23222_1080# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X494 XA20.XA1.MP0.S SARP XA20.XA1.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X495 XA6.XA9.MN1.S XA6.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R56 XDAC1.XC128b<2>.XRES1B.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X496 AVSS XA0.CMP_OP XA4.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X497 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X498 XA6.CN0 XA6.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X499 AVSS XA4.CN1 D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R57 XDAC1.X16ab.XRES16.B XA2.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X500 VREF XA2.XA2.A XA2.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R58 XDAC1.XC0.XRES2.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X501 D<2> XA6.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X502 XA4.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X503 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X504 AVDD XA0.XA6.Y XA0.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X505 XA2.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X506 XA6.XA1.XA4.MN2.S XA6.XA1.XA4.LCK_N XA6.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X507 XA2.DONE XA2.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X508 XA5.CP0 XA5.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X509 XA5.CP0 XA5.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X510 D<5> XA3.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X511 D<5> XA3.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R59 XA1.CN0 XDAC2.XC64a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X512 XA0.CP1 D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X513 XA5.CN1 XA5.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X514 XA2.CN0 XA2.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X515 XA5.CN1 XA5.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X516 AVSS XA6.XA2.A XA6.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X517 XA2.CEO XA2.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X518 XA5.ENO XA5.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X519 AVDD XA5.XA1.XA1.MP3.G XA5.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X520 XA20.XA3.N2 SARN XA20.XA2.N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X521 XA20.XA2.VMR XA20.XA1.CK AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R60 XB2.XA4.GNG m3_23222_120# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X522 XA2.XA8.A XA2.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X523 XA8.XA1.CHL_OP XA7.ENO XA8.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X524 XB2.CKN CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R61 XDAC1.XC64b<1>.XRES8.B D<7> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X525 VREF XA2.XA1.CHL_OP XA2.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X526 XA20.XA4.MP0.S SARN XA20.XA4.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X527 D<1> XA7.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X528 D<1> XA7.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X529 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X530 XA6.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X531 XA4.XA1.CHL_OP EN XA4.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X532 XA5.CN1 XA5.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X533 VREF XA8.XA2.A XA8.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X534 AVSS XA0.CEO XA1.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X535 XA5.CN1 XA5.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X536 XA3.XA1.XA5.MN2.S XA3.XA1.XA4.LCK_N XA3.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X537 XA1.XA11.Y XA0.CEO XA1.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X538 XA3.XA1.XA5.MP2.S EN XA3.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R62 XA1.CN0 XDAC2.XC64a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X539 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X540 XA0.XA1.XA5.MN2.S XA0.XA1.XA4.LCK_N XA0.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X541 XA5.XA1.XA4.LCK_N XA5.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X542 XA8.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X543 XA1.XA6.Y CK_SAMPLE XA1.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X544 XA5.XA1.XA4.LCK_N XA5.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X545 XA1.XA6.Y D<7> XA1.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X546 DONE XA8.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 AVSS XA1.XA1.CHL_OP XA1.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X548 VREF XA1.XA1.CHL_OP XA1.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R63 XDAC1.XC32a<0>.XRES8.B D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R64 XDAC1.XC1.XRES1B.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X549 XA6.XA1.XA1.MN2.S XA5.ENO XA6.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X550 XA4.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 XA8.CN0 XA8.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X552 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X553 XA4.XA9.MN1.S XA4.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R65 XDAC1.XC64a<0>.XRES16.B XA1.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X554 XA8.CEO XA8.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X555 AVSS CK_SAMPLE XA1.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R66 XA0.CN0 XDAC2.XC128b<2>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X556 XA7.XA1.XA5.MN2.S XA7.XA1.XA4.LCK_N XA7.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X557 AVDD XA1.CN0 XA1.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X558 XA4.CN0 XA4.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X559 XA7.XA1.XA5.MP2.S EN XA7.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X560 XA8.XA8.A XA8.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X561 VREF XA0.XA2.A D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X562 D<4> XA4.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X563 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R67 XDAC1.X16ab.XRES8.B XA3.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X564 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X565 VREF XA8.XA1.CHL_OP XA8.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X566 XB1.XA1.MP0.G XB1.XA1.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X567 XA4.XA1.XA4.MN2.S XA4.XA1.XA4.LCK_N XA4.XA1.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X568 XA0.DONE XA0.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X569 XA0.CN0 XA0.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X570 XA6.CP0 XA6.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X571 AVSS XA4.XA2.A XA4.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X572 XA0.CEO XA0.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R68 D<8> XDAC2.XC128a<1>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X573 XA6.CN1 XA6.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R69 XDAC1.XC64a<0>.XRES8.B XA1.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X574 XA2.XA11.MP1.S XA2.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X575 XA0.XA8.A XA0.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X576 XA6.XA11.Y XA5.CEO XA6.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X577 XA6.ENO XA6.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X578 XA2.XA6.MP3.S D<6> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X579 VREF XA0.XA1.CHL_OP XA0.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X580 D<3> XA5.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X581 D<3> XA5.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R70 XDAC1.X16ab.XRES1A.B D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X582 XA4.XA1.XA1.MN2.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X583 XA6.XA6.Y D<2> XA6.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X584 XA2.CP0 XA2.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X585 XA20.XA4.MP0.S SARN XA20.XA4.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X586 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X587 VREF XA6.XA1.CHL_OP XA6.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X588 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X589 XA2.XA10.Y XA2.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X590 AVSS XB1.CKN XB1.XA3.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X591 XA2.XA2.A EN XA2.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R71 D<8> XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X592 XA3.XA1.CHL_OP XA2.ENO XA3.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X593 AVSS XA20.XA2.CO XA0.CMP_ON AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X594 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X595 XA3.XA1.CHL_OP EN XA3.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X596 AVDD XA20.XA2.CO XA0.CMP_ON AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X597 XA6.CN1 XA6.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X598 XA0.XA1.CHL_OP EN XA0.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X599 AVSS XA1.CEO XA2.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X600 XA2.XA6.MP1.S XA2.CN0 XA2.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X601 XA2.XA1.XA1.MP3.S XA0.CMP_OP XA2.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R72 m3_16526_1240# XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X602 XA4.XA1.XA1.MN2.S XA4.EN XA4.XA1.XA1.MP3.G AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X603 AVDD XA6.CN0 XA6.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X604 XA2.XA6.Y CK_SAMPLE XA2.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R73 D<8> XDAC2.XC128a<1>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X605 XA6.XA1.XA4.LCK_N XA6.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X606 VREF XA2.CN1 D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X607 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X608 AVDD XA20.XA1.CKN XA20.XA4.MP0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X609 XA20.XA4.MP0.S XA20.XA1.CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X610 AVSS XA2.XA1.CHL_OP XA2.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X611 XA2.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X612 XA5.XA1.XA5.MN2.S XA5.XA1.XA4.LCK_N XA5.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X613 SAR_IP XB1.M1.G SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X614 XA5.XA1.XA5.MP2.S EN XA5.XA1.XA5.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X615 XA3.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R74 XDAC1.XC128b<2>.XRES16.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X616 XA3.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X617 XA8.XA11.MP1.S XA8.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X618 XA0.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R75 XA0.CN0 XDAC2.XC128b<2>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X619 SAR_IN XB1.TIE_L SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X620 AVSS XA1.CP0 XA1.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X621 XA7.XA1.CHL_OP XA6.ENO XA7.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X622 XA7.XA1.CHL_OP EN XA7.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X623 VREF XA1.CP0 XA1.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X624 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X625 AVSS CK_SAMPLE XA2.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X626 XA8.XA6.MP3.S D<0> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R76 XA1.CN1 XDAC2.XC64b<1>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X627 AVSS XA1.CN1 D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X628 XA20.XA10.A DONE XA20.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X629 AVSS DONE XA20.XA10.A AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X630 VREF XA1.CN1 D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X631 XA8.CP0 XA8.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X632 XB1.XA4.MN1.S XB1.CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X633 XA8.XA10.Y XA8.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X634 AVSS XA1.CP0 XA1.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X635 SAR_IN XB1.TIE_L SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X636 XA7.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X637 XA8.XA2.A EN XA8.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X638 VREF XA1.CP0 XA1.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X639 XA4.CP0 XA4.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X640 XA7.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X641 AVSS XA7.CEO XA8.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X642 XA8.XA6.MP1.S XA8.CN0 XA8.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R77 XA1.CN0 XDAC2.XC64a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X643 SAR_IN XB2.M1.G SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R78 m3_830_3960# XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X644 XA8.XA1.XA1.MP3.S XA0.CMP_OP XA8.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X645 XA4.CN1 XA4.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X646 XA0.XA11.MP1.S XA0.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R79 AVSS XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X647 XA8.XA6.Y CK_SAMPLE XA8.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X648 VREF XA8.CN1 D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X649 XA20.XA1.MP0.S SARP XA20.XA1.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
R80 D<8> XDAC2.XC128a<1>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X650 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X651 XA4.XA11.Y XA4.CEIN XA4.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X652 XA4.ENO XA4.XA1.XA1.MP3.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X653 XA0.XA6.MP3.S XA0.CP1 AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X654 XA1.XA10.A XA1.XA6.Y XA1.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X655 AVSS XA8.XA1.CHL_OP XA8.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X656 XA8.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X657 AVDD XA1.XA6.Y XA1.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X658 XA4.XA6.Y D<4> XA4.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X659 XA0.CP0 XA0.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X660 VREF XA4.XA1.CHL_OP XA4.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X661 D<2> XA6.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X662 XA0.XA10.Y XA0.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X663 AVSS CK_SAMPLE XA8.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X664 XA0.XA2.A EN XA0.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R81 m3_830_120# XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
R82 XA1.CN1 XDAC2.XC64b<1>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X665 XA4.CN1 XA4.XA2.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R83 XB1.XA3.B m3_7598_3160# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
R84 D<8> XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X666 XA2.XA10.A XA2.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X667 XA0.XA6.MP1.S XA0.CN0 XA0.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X668 XA0.XA1.XA1.MP3.S XA0.CMP_OP XA0.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X669 AVDD XA4.CN0 XA4.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X670 XA4.XA1.XA4.LCK_N XA4.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X671 XA2.CN0 XA2.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X672 VREF D<8> XA0.CP1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X673 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X674 VREF XA6.CP0 XA6.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X675 XA0.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R85 D<8> XDAC2.XC128a<1>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X676 D<6> XA2.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X677 VREF XA6.CN1 D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R86 XDAC1.XC1.XRES1A.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R87 XA7.CN0 XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X678 XA5.XA1.CHL_OP XA4.ENO XA5.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X679 XA2.XA1.XA4.MP2.S EN XA2.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X680 AVSS XA20.XA2.VMR XA0.CMP_OP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X681 AVDD XB2.CKN XB2.XA3.MP0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X682 XA5.XA1.CHL_OP EN XA5.XA1.XA4.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X683 AVDD XA20.XA2.VMR XA0.CMP_OP AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X684 XA6.XA1.XA5.MN2.S XA6.XA1.XA4.LCK_N XA6.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X685 XB2.CKN CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X686 VREF XA6.CP0 XA6.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R88 XDAC1.XC64a<0>.XRES1B.B XA1.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R89 XA3.CN1 XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R90 XA1.CN1 XDAC2.XC64b<1>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X687 AVSS XA2.CP0 XA2.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X688 VREF XA2.XA2.A XA2.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X689 XA20.XA1.CKN XA20.XA10.B XA20.XA10.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X690 AVDD XA20.XA10.B XA20.XA1.CKN AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X691 AVSS XA2.CN1 D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X692 XA5.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X693 XA5.XA1.XA4.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X694 XA8.XA10.A XA8.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X695 AVDD XA6.XA6.Y XA6.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X696 AVSS XA2.CP0 XA2.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X697 XA8.CN0 XA8.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X698 XB1.TIE_L XB1.XA2.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X699 XA2.XA1.XA1.MP2.S XA0.CMP_ON XA2.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X700 AVSS XA1.XA2.A XA1.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X701 VREF XA1.XA2.A XA1.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R91 XA0.CN0 XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R92 XB1.XA3.B m3_7598_280# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
R93 XA6.CN0 XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X702 D<0> XA8.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X703 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X704 XA20.XA3.N2 SARN XA20.XA2.N1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X705 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X706 XA20.XA2.VMR XA20.XA2.CO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X707 AVSS XA2.CEO XA3.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X708 XA8.XA1.XA4.MP2.S EN XA8.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X709 XA3.XA11.Y XA2.CEO XA3.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X710 XA1.DONE XA1.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X711 AVSS XB1.TIE_L XA0.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X712 XA1.DONE XA1.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X713 D<4> XA4.CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X714 AVDD EN XA2.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X715 XA2.XA10.A XA2.XA6.Y XA2.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X716 XA3.XA6.Y CK_SAMPLE XA3.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X717 XA3.XA6.Y D<5> XA3.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X718 XA1.CN0 XA1.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X719 XA1.CN0 XA1.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X720 XA0.XA10.A XA0.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X721 XA0.XA6.Y CK_SAMPLE XA0.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X722 AVSS XA8.CP0 XA8.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X723 VREF XA8.XA2.A XA8.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X724 XA1.CEO XA1.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X725 AVSS XA3.XA1.CHL_OP XA3.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X726 XA1.CEO XA1.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X727 AVSS XA0.XA1.CHL_OP XA0.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X728 VREF XA3.XA1.CHL_OP XA3.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R94 D<8> XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X729 XA0.CN0 XA0.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X730 XA1.XA8.A XA1.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X731 AVSS XA8.CN1 D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X732 XB1.XA3.B XB1.CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X733 XA1.XA8.A XA1.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R95 XDAC1.XC128b<2>.XRES2.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X734 VREF XA4.CP0 XA4.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X735 AVSS XA6.CEO XA7.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X736 XA0.CP1 D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X737 XA7.XA11.Y XA6.CEO XA7.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X738 AVSS CK_SAMPLE XA3.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X739 AVSS XA1.XA1.CHL_OP XA1.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X740 AVSS CK_SAMPLE XA0.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X741 AVDD XA3.CN0 XA3.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X742 VREF XA1.XA1.CHL_OP XA1.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X743 VREF XA4.CN1 D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X744 AVSS XA8.CP0 XA8.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R96 m3_16526_4120# XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X745 XA8.XA1.XA1.MP2.S XA0.CMP_ON XA8.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X746 XA7.XA6.Y CK_SAMPLE XA7.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X747 XA0.XA1.XA4.MP2.S EN XA0.XA1.XA4.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X748 XA7.XA6.Y D<1> XA7.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X749 XA4.XA1.XA5.MN2.S XA4.XA1.XA4.LCK_N XA4.XA1.XA5.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X750 AVSS XA7.XA1.CHL_OP XA7.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X751 SAR_IP XB1.TIE_L SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X752 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X753 VREF XA4.CP0 XA4.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X754 VREF XA7.XA1.CHL_OP XA7.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X755 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X756 AVDD XB2.M1.G XB2.XA4.GNG AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X757 XA6.XA1.CHL_OP XA5.ENO XA6.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X758 XA2.CP0 XA2.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X759 VREF XA0.XA2.A D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R97 XA3.CN1 XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R98 XA1.CN1 XDAC2.XC64b<1>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X760 AVDD EN XA8.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X761 XA8.XA10.A XA8.XA6.Y XA8.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X762 AVSS CK_SAMPLE XA7.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X763 XA2.CN1 XA2.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X764 AVDD XA7.CN0 XA7.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X765 XB2.M1.G XB2.XA1.Y XB2.XA4.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X766 VREF XA6.XA2.A XA6.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R99 XDAC1.XC128a<1>.XRES8.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R100 D<8> XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X767 SAR_IP XB1.TIE_L SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X768 AVDD XA2.XA1.XA1.MP3.G XA2.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X769 AVDD XA4.XA6.Y XA4.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R101 m3_830_3000# XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X770 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X771 XA0.XA1.XA1.MP2.S XA0.CMP_ON XA0.ENO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X772 XA6.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X773 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X774 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X775 XA6.DONE XA6.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X776 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X777 AVDD XA20.XA1.CK XA20.XA4.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X778 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X779 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X780 XA6.CN0 XA6.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X781 AVSS XA2.XA2.A XA2.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X782 XA2.CN1 XA2.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X783 XA20.XA2.N1 SARN XA20.XA3.N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R102 XDAC1.XC0.XRES4.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X784 AVDD EN XA0.XA1.XA1.MP3.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X785 XA6.CEO XA6.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X786 AVDD AVDD XA20.XA3.N2 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R103 XA0.CN0 XDAC2.XC128b<2>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X787 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X788 XA20.XA10.B XA8.CEO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X789 XA2.XA1.XA4.LCK_N XA2.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X790 XA20.XA10.B XA8.CEO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X791 XA6.XA8.A XA6.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R104 XB2.XA4.GNG m3_23222_2040# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X792 XA0.CMP_OP XA20.XA2.VMR AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X793 XA8.CP0 XA8.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X794 XA0.CMP_OP XA20.XA2.VMR AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X795 XA2.DONE XA2.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R105 XDAC1.XC128a<1>.XRES1A.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R106 XDAC1.XC1.XRES2.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X796 XA20.XA4.MP0.S SARN XA20.XA4.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X797 XA20.XA1.MP0.S SARP XA20.XA1.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X798 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X799 VREF XA6.XA1.CHL_OP XA6.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X800 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X801 XA2.CN0 XA2.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X802 XA8.CN1 XA8.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X803 XA1.XA11.Y XA1.XA10.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X804 XA20.XA2.N1 XA20.XA1.CK AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X805 XA1.XA11.MP1.S XA1.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 AVDD XA20.XA1.CK XA20.XA2.N1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X807 XA2.CEO XA2.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X808 AVSS XA4.CEO XA5.XA11.Y AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X809 XA5.XA11.Y XA4.CEO XA5.XA11.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X810 AVDD XA8.XA1.XA1.MP3.G XA8.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X811 XA1.XA6.MN3.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R107 XDAC1.XC128b<2>.XRES4.B XA0.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X812 XA20.XA2.CO XA20.XA2.VMR XA20.XA2.N2 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X813 XA1.XA6.MP3.S D<7> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X814 AVDD XA20.XA2.VMR XA20.XA2.CO AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X815 XA2.XA8.A XA2.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X816 XA5.XA6.Y CK_SAMPLE XA5.XA6.MN3.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X817 XA5.XA6.Y D<3> XA5.XA6.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X818 AVSS XA3.CP0 XA3.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R108 XDAC1.XC64b<1>.XRES1A.B D<7> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X819 SAR_IN XB2.M1.G SARN AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X820 VREF XA3.CP0 XA3.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X821 XA1.CP0 XA1.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X822 XA1.CP0 XA1.XA1.CHL_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X823 AVSS XA0.CP0 XA0.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X824 AVSS XA2.XA1.CHL_OP XA2.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X825 AVSS XA5.XA1.CHL_OP XA5.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X826 XA1.XA10.Y XA1.XA10.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X827 VREF XA5.XA1.CHL_OP XA5.CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X828 AVSS XA3.CN1 D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X829 XA1.XA2.A XA0.ENO XA1.XA1.XA5.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R109 XA0.CN0 XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X830 XA1.XA10.Y XA1.XA10.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X831 AVSS D<8> XA0.CP1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X832 VREF XA3.CN1 D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X833 XA1.XA2.A EN XA1.XA1.XA5.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X834 XA0.CP0 XA0.XA1.CHL_OP VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X835 XA4.XA1.CHL_OP XA4.EN XA4.XA1.XA4.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X836 XA1.XA6.MN1.S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X837 XA8.CN1 XA8.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X838 AVSS XA8.XA2.A XA8.CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X839 SAR_IP XB1.M1.G SARP AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X840 XA1.XA6.MP1.S XA1.CN0 XA1.XA6.Y AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X841 AVSS XA0.CMP_OP XA1.XA1.XA1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X842 XA1.XA1.XA1.MP3.S XA0.CMP_OP XA1.XA1.XA1.MP2.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X843 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X844 AVSS CK_SAMPLE XA5.XA6.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X845 D<8> XA0.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X846 AVDD XB1.M1.G XB1.XA4.GNG AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X847 AVDD XA5.CN0 XA5.XA6.MP1.S AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X848 AVSS XA3.CP0 XA3.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X849 AVSS XA1.CN1 D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R110 XDAC1.XC64a<0>.XRES4.B XA1.CP0 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X850 XA8.XA1.XA4.LCK_N XA8.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X851 AVSS XA0.CP0 XA0.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X852 VREF XA3.CP0 XA3.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X853 VREF XA1.CN1 D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X854 VREF XA4.XA2.A XA4.CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X855 DONE XA8.XA8.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X856 AVSS XA7.CP0 XA7.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X857 AVDD XA0.XA1.XA1.MP3.G XA0.XA1.XA1.MP3.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X858 VREF XA7.CP0 XA7.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X859 XA1.XA1.XA5.MN1.S XA0.CMP_ON AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R111 XDAC1.XC32a<0>.XRES1A.B AVSS sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X860 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X861 XA1.XA1.XA5.MP1.S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R112 XDAC1.XC128a<1>.XRES1B.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R113 XB1.XA3.B m3_7598_1240# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X862 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X863 XA4.XA1.XA4.MN1.S XA0.CMP_OP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X864 XA8.CN0 XA8.CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X865 AVSS XA7.CN1 D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X866 VREF XA7.CN1 D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X867 XA4.DONE XA4.XA8.A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X868 XA8.CEO XA8.XA11.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X869 D<6> XA2.CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X870 XA3.XA10.A XA3.XA6.Y XA3.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X871 XA0.XA10.A XA0.XA6.Y XA0.XA9.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X872 AVDD XA3.XA6.Y XA3.XA10.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X873 XA4.CN0 XA4.CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X874 XA8.XA8.A XA8.ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X875 AVSS XA7.CP0 XA7.CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X876 D<8> XA0.XA2.A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X877 VREF XA7.CP0 XA7.CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X878 XA4.CEO XA4.XA11.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R114 XDAC1.XC64b<1>.XRES1B.B D<7> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X879 AVSS XA8.XA1.CHL_OP XA8.CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X880 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R115 XDAC1.XC0.XRES16.B XA0.CP1 sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X881 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X882 AVSS XB2.CKN XB2.XA3.MP0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X883 XA0.XA1.XA4.LCK_N XA0.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X884 XA4.XA8.A XA4.ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X885 XA6.XA11.MP1.S XA6.XA10.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 XA2.XA1.CHL_OP a_4862_42588# 0.01727f
C1 XA7.XA1.CHL_OP XA0.CMP_OP 0.03343f
C2 XA0.XA10.A AVDD 0.769273f
C3 XA0.CMP_OP a_13574_40828# 0.014652f
C4 XA1.XA1.XA4.LCK_N a_2342_41180# 0.023475f
C5 XA20.XA10.B XA20.XA11.MP1.S 0.026506f
C6 XA6.XA1.XA1.MP3.S a_16094_40476# 0.04865f
C7 a_9902_46108# CK_SAMPLE 0.073189f
C8 a_12422_46108# AVDD 0.378183f
C9 XA8.XA6.MP1.S VREF 0.011406f
C10 XA20.XA4.MP0.S SARN 0.253395f
C11 a_4862_49804# a_4862_49452# 0.010937f
C12 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES2.B 0.015267f
C13 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES8.B 0.477132f
C14 a_21134_45228# XA8.XA1.CHL_OP 0.066018f
C15 XA7.ENO XA7.XA1.XA4.LCK_N 0.154232f
C16 XB2.XA4.GNG m3_23150_3000# 0.024512f
C17 XB1.XA3.B m3_830_120# 0.172147f
C18 XA4.CEIN AVDD 1.04893f
C19 a_13574_48572# a_13574_48220# 0.010937f
C20 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES1A.B 0.022835f
C21 XDAC1.XC64a<0>.XRES8.B XDAC1.XC64a<0>.XRES16.B 0.1057f
C22 XA4.XA1.XA5.MN2.S XA4.XA1.XA5.MN1.S 0.050207f
C23 a_4862_46988# CK_SAMPLE 0.070402f
C24 XA6.ENO VREF 0.879117f
C25 XA8.ENO D<0> 0.402335f
C26 a_7382_46988# AVDD 0.395571f
C27 XA4.ENO EN 1.02916f
C28 XA0.XA1.XA4.LCK_N D<8> 0.033627f
C29 XA0.XA1.XA5.MN2.S EN 0.027112f
C30 XA2.ENO XA2.XA2.A 0.090222f
C31 a_16094_39772# AVDD 0.382569f
C32 XA0.XA10.Y a_974_48572# 0.091063f
C33 XA5.XA11.MP1.S XA5.XA10.Y 0.010335f
C34 XA4.EN XA3.XA1.XA1.MP2.S 0.155821f
C35 XA2.ENO XA3.XA1.XA1.MN2.S 0.038148f
C36 XA6.XA2.A a_14942_42588# 0.089492f
C37 XA0.XA2.A XA0.XA1.XA5.MN2.S 0.050207f
C38 XDAC1.XC128b<2>.XRES8.B SARP 27.705599f
C39 XA0.CMP_OP a_7382_40124# 0.066394f
C40 XA8.XA6.Y AVDD 0.860513f
C41 XA0.XA6.Y XA0.ENO 0.051732f
C42 XA4.XA6.Y VREF 0.078171f
C43 XA5.XA1.XA1.MN2.S a_13574_40124# 0.056787f
C44 XA6.XA8.A a_14942_47692# 0.160931f
C45 XA0.XA8.A a_974_47340# 0.091063f
C46 XA3.XA6.Y XA3.DONE 0.014904f
C47 XA3.CN1 AVDD 2.00341f
C48 XB2.XA1.MP0.G XB2.CKN 0.015687f
C49 a_12422_2094# a_12422_1742# 0.010937f
C50 a_13862_1918# XB2.M1.G 0.036098f
C51 XB1.M1.G XB1.XA4.GNG 0.250687f
C52 XA7.XA1.XA1.MP3.S AVDD 0.139093f
C53 XA1.CEO a_4862_49100# 0.070731f
C54 XA1.XA11.Y a_3494_49100# 0.104051f
C55 a_14942_49452# a_14942_49100# 0.010937f
C56 XDAC1.X16ab.XRES16.B XDAC1.X16ab.XRES1A.B 0.467299f
C57 XA2.CN1 a_6014_43468# 0.070763f
C58 XA6.XA1.CHL_OP XA0.CMP_OP 0.033149f
C59 XA4.ENO a_11054_41180# 0.072087f
C60 XDAC2.XC0.XRES2.B SARN 7.01089f
C61 a_13574_48220# XA5.XA6.Y 0.071154f
C62 XA6.XA1.XA1.MP3.G a_16094_40476# 0.098305f
C63 a_8534_46108# CK_SAMPLE 0.07476f
C64 a_6014_46108# D<6> 0.011483f
C65 a_11054_46108# AVDD 0.378183f
C66 XA7.XA6.Y XA7.CP0 0.010942f
C67 XA2.ENO XA2.CN0 0.093196f
C68 XA0.XA1.XA4.MP1.S EN 0.027563f
C69 XA5.XA1.XA4.MP2.S AVDD 0.035519f
C70 a_19982_45228# XA8.XA1.CHL_OP 0.06825f
C71 XA6.ENO XA7.XA1.XA4.LCK_N 0.3401f
C72 XA7.ENO XA8.XA1.XA5.MN2.S 0.010423f
C73 XB2.XA4.GNG m3_16598_3160# 0.0666f
C74 XB1.XA3.B m3_7598_280# 0.024512f
C75 a_11054_2798# SAR_IP 0.02841f
C76 a_12422_2798# SARP 0.010335f
C77 XA2.XA11.Y AVDD 0.712901f
C78 XA0.XA10.A a_974_48220# 0.070424f
C79 a_18614_41180# a_18614_40828# 0.010937f
C80 XA0.CN0 XDAC2.XC128b<2>.XRES16.B 0.028741f
C81 a_3494_46988# CK_SAMPLE 0.068905f
C82 XA5.ENO VREF 0.879117f
C83 a_2342_46988# D<7> 0.070283f
C84 a_6014_46988# AVDD 0.395571f
C85 XA4.EN EN 0.952619f
C86 a_12422_39772# a_12422_39420# 0.010937f
C87 XA2.XA6.Y XA2.XA6.MP1.S 0.055045f
C88 XA3.XA1.XA5.MP2.S AVDD 0.038567f
C89 a_21134_42588# EN 0.077363f
C90 a_13862_334# a_13862_n18# 0.010937f
C91 a_11054_46108# XA4.CP0 0.066018f
C92 XA1.ENO XA2.XA2.A 0.04064f
C93 XA0.CP1 XA3.CN1 0.145077f
C94 XA0.XA10.Y a_n178_48572# 0.13253f
C95 XA3.XA1.CHL_OP a_8534_41884# 0.040867f
C96 XA0.CMP_ON XA3.XA1.XA4.LCK_N 0.284482f
C97 XA0.CMP_ON a_21134_39772# 0.067588f
C98 XA6.XA1.XA4.MN2.S XA6.XA1.XA4.MN1.S 0.050207f
C99 XA0.CMP_OP a_6014_40124# 0.067964f
C100 XA7.XA6.Y CK_SAMPLE 0.179573f
C101 XA0.XA8.A a_n178_47340# 0.127528f
C102 XA2.CN1 AVDD 2.00391f
C103 XB1.M1.G XB2.M1.G 0.017476f
C104 XA20.XA1.CKN XA20.XA2.N1 0.038766f
C105 XB1.TIE_L a_13862_2974# 0.03839f
C106 XA3.CN0 XA7.CN0 0.071907f
C107 XA4.XA1.XA1.MP3.G D<4> 0.021797f
C108 XA0.XA1.XA1.MP3.G EN 0.176792f
C109 XA7.XA1.XA1.MP3.G AVDD 1.05472f
C110 a_23654_40828# SARP 0.023578f
C111 XA5.CEO XA6.XA11.Y 0.220689f
C112 XA1.XA11.Y a_2342_49100# 0.089492f
C113 XA2.CN1 a_4862_43468# 0.111278f
C114 XA1.XA1.CHL_OP a_3494_42588# 0.01727f
C115 XA8.XA1.CHL_OP XA8.XA2.A 0.133602f
C116 XA5.XA1.CHL_OP XA0.CMP_OP 0.03343f
C117 XA4.ENO a_9902_41180# 0.068502f
C118 XDAC1.XC0.XRES8.B SARP 27.705502f
C119 a_22502_48572# AVDD 0.471468f
C120 XDAC2.XC32a<0>.XRES16.B SARN 55.2956f
C121 XA8.XA10.A XA8.XA8.A 0.062692f
C122 a_12422_48220# XA5.XA6.Y 0.067588f
C123 XA6.XA1.XA1.MP3.G a_14942_40476# 0.066018f
C124 XA1.XA1.XA1.MP3.G XA1.XA1.XA1.MN2.S 0.078539f
C125 XA1.XA1.XA1.MP3.S XA1.XA1.XA1.MP2.S 0.050207f
C126 XA8.CN0 VREF 0.452875f
C127 XA8.XA6.MP1.S D<0> 0.016737f
C128 XA4.XA1.XA4.MP2.S AVDD 0.035519f
C129 a_3494_49804# a_3494_49452# 0.010937f
C130 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES8.B 0.477132f
C131 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES2.B 0.015267f
C132 XA1.XA1.CHL_OP XA2.XA1.CHL_OP 0.082663f
C133 XA3.CP0 XA3.CN1 0.183039f
C134 XB2.XA1.MP0.G AVDD 0.518987f
C135 XB2.XA4.GNG m3_16526_3160# 0.105547f
C136 XB1.XA3.B m3_7526_280# 0.024512f
C137 XA2.CEO AVDD 1.98375f
C138 a_12422_48572# a_12422_48220# 0.010937f
C139 XA0.XA10.A a_n178_48220# 0.132671f
C140 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES16.B 0.063821f
C141 XDAC2.XC64a<0>.XRES8.B XDAC2.XC64a<0>.XRES2.B 0.446669f
C142 XA7.ENO D<1> 0.499068f
C143 XA4.ENO VREF 0.879117f
C144 XA2.ENO EN 1.02916f
C145 XA8.XA6.Y a_21134_46988# 0.023982f
C146 XA3.XA6.Y XA3.XA6.MN3.S 0.089305f
C147 XA2.XA6.Y XA2.XA6.MN1.S 0.026506f
C148 XA2.XA1.XA5.MP2.S AVDD 0.038567f
C149 XA0.CP1 XA2.CN1 0.147379f
C150 XA4.CN0 XA4.XA1.CHL_OP 0.037542f
C151 a_9902_46108# XA4.CP0 0.067789f
C152 XA1.ENO XA1.XA2.A 0.090222f
C153 XA2.ENO XA2.XA1.XA1.MP2.S 0.150467f
C154 XA20.XA2.N1 a_23654_42236# 0.031884f
C155 XA3.XA1.CHL_OP a_7382_41884# 0.023777f
C156 XA5.XA2.A a_13574_42588# 0.091063f
C157 XA0.CMP_ON a_19982_39772# 0.066018f
C158 XA0.CMP_OP a_4862_40124# 0.072221f
C159 XA5.XA6.Y D<3> 0.039903f
C160 XA3.XA8.A VREF 0.028938f
C161 XA7.XA8.A AVDD 1.19556f
C162 XA5.XA1.XA1.MP3.G a_13574_39420# 0.023111f
C163 XA5.XA1.XA1.MP2.S a_12422_40124# 0.04865f
C164 XA1.CN1 AVDD 2.00341f
C165 XA6.XA6.Y a_14942_47692# 0.017683f
C166 a_7382_44348# VREF 0.059568f
C167 XA2.XA8.A XA2.DONE 0.1303f
C168 a_11054_2094# a_11054_1742# 0.010937f
C169 a_8462_1918# XB1.XA4.GNG 0.01152f
C170 XA0.XA1.XA1.MP3.G D<8> 0.012174f
C171 XA6.XA1.XA1.MP3.S AVDD 0.139596f
C172 a_13574_49452# a_13574_49100# 0.010937f
C173 XA5.CEO XA6.CEO 0.033943f
C174 XDAC2.X16ab.XRES2.B XDAC2.X16ab.XRES1A.B 0.015267f
C175 XA4.XA1.CHL_OP XA0.CMP_OP 0.033149f
C176 a_21134_48572# AVDD 0.394716f
C177 XDAC1.XC32a<0>.XRES2.B SARP 7.01089f
C178 XA0.CMP_OP a_9902_40828# 0.014592f
C179 XA8.XA10.A XA8.XA9.MN1.S 0.073313f
C180 XA20.XA10.B XA20.XA10.A 0.412143f
C181 XA1.XA1.XA1.MP3.G XA1.XA1.XA1.MP2.S 0.064105f
C182 XA1.XA1.XA4.MP2.S EN 0.027192f
C183 XA6.CN0 XA6.XA2.A 0.035589f
C184 a_18614_45228# XA7.XA1.CHL_OP 0.066679f
C185 XA2.CP0 XA3.CN1 0.135532f
C186 XA3.CP0 XA2.CN1 0.065837f
C187 XA6.ENO XA7.XA1.XA5.MN2.S 0.010423f
C188 a_15014_2270# AVDD 0.470727f
C189 XB2.XA4.GNG m3_23222_3960# 0.049023f
C190 XB1.XA3.B m3_974_1080# 0.0666f
C191 XA1.XA11.Y AVDD 0.708074f
C192 XA3.XA1.XA4.LCK_N XA3.XA1.XA5.MN1.S 0.030434f
C193 XA4.XA1.XA5.MN2.S XA4.XA1.XA4.LCK_N 0.010898f
C194 XA7.ENO a_19982_39420# 0.071936f
C195 a_17462_41180# a_17462_40828# 0.010937f
C196 XA6.ENO D<1> 0.071215f
C197 XA4.EN VREF 0.879117f
C198 XA1.ENO EN 0.952619f
C199 a_11054_39772# a_11054_39420# 0.010937f
C200 XA8.XA6.Y a_19982_46988# 0.047651f
C201 a_21134_42588# VREF 0.028416f
C202 XA2.XA1.XA4.LCK_N AVDD 0.271451f
C203 XA1.XA1.XA4.LCK_N D<7> 0.01587f
C204 XA2.XA6.Y XA2.CN0 0.093605f
C205 a_12422_334# a_12422_n18# 0.010937f
C206 XA0.CP1 XA1.CN1 1.77286f
C207 XA0.ENO XA1.XA2.A 0.041437f
C208 a_12422_39772# AVDD 0.382762f
C209 XA5.CEO XA5.XA10.A 0.010854f
C210 XA8.CEO a_23654_48572# 0.066372f
C211 XDAC2.XC128a<1>.XRES1A.B XDAC2.XC32a<0>.XRES1B.B 0.62895f
C212 XA2.ENO XA2.XA1.XA1.MN2.S 0.040976f
C213 XA8.ENO a_21134_40476# 0.017019f
C214 XA5.XA2.A a_12422_42588# 0.127528f
C215 XDAC2.XC128b<2>.XRES8.B SARN 27.705599f
C216 XA0.CMP_ON a_18614_39772# 0.067588f
C217 XA0.CMP_OP a_3494_40124# 0.073806f
C218 XA3.XA6.Y VREF 0.078171f
C219 XA7.XA6.Y AVDD 0.864413f
C220 XA5.XA1.XA1.MP3.G a_12422_39420# 0.03422f
C221 a_21134_44348# AVDD 0.377363f
C222 a_6014_44348# VREF 0.059568f
C223 a_12422_44348# D<3> 0.02026f
C224 XA0.CN0 a_974_46108# 0.103403f
C225 XA6.XA1.XA1.MP3.G AVDD 1.07016f
C226 XA0.CEO a_3494_49100# 0.0733f
C227 XA5.CEO XA5.XA11.Y 0.377598f
C228 XA1.CN1 a_3494_43468# 0.112954f
C229 XA7.XA1.CHL_OP XA7.XA2.A 0.133602f
C230 XA3.XA1.CHL_OP XA0.CMP_OP 0.03343f
C231 XA4.EN a_8534_41180# 0.06753f
C232 XA0.CMP_OP a_8534_40828# 0.014652f
C233 XA0.XA9.MN1.S XA0.XA8.A 0.010335f
C234 a_4862_46108# CK_SAMPLE 0.073189f
C235 XA8.CN0 D<0> 0.437663f
C236 a_7382_46108# AVDD 0.378183f
C237 XA0.XA1.XA4.MP2.S EN 0.027664f
C238 XA3.XA1.XA4.MP1.S AVDD 0.105303f
C239 a_2342_49804# a_2342_49452# 0.010937f
C240 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES8.B 0.029725f
C241 XDAC2.XC0.XRES16.B XDAC2.XC64b<1>.XRES16.B 0.010386f
C242 a_17462_45228# XA7.XA1.CHL_OP 0.067588f
C243 XA2.CP0 XA2.CN1 0.114645f
C244 XA1.CP0 XA3.CN1 0.13878f
C245 XA3.CP0 XA1.CN1 0.071833f
C246 XB1.XA3.B m3_830_1080# 0.172147f
C247 XB2.XA4.GNG m3_23150_3960# 0.024512f
C248 XA1.CEO AVDD 1.04893f
C249 a_23654_48572# XA20.XA10.B 0.023111f
C250 a_11054_48572# a_11054_48220# 0.010937f
C251 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES16.B 0.063821f
C252 XDAC1.XC64a<0>.XRES8.B XDAC1.XC64a<0>.XRES2.B 0.446669f
C253 a_n178_46988# CK_SAMPLE 0.070402f
C254 XA2.ENO VREF 0.879117f
C255 XA6.ENO D<2> 0.431648f
C256 a_2342_46988# AVDD 0.395571f
C257 XA0.ENO EN 1.04628f
C258 a_17462_42588# EN 0.078934f
C259 a_8534_46108# XA3.CP0 0.066219f
C260 XA0.ENO XA0.XA2.A 0.090222f
C261 a_11054_39772# AVDD 0.382569f
C262 XA8.CEO a_22502_48572# 0.077615f
C263 XA4.XA10.Y XA4.XA11.MP1.S 0.010335f
C264 XA2.XA1.CHL_OP a_6014_41884# 0.023777f
C265 XA1.ENO XA2.XA1.XA1.MN2.S 0.030034f
C266 XDAC1.XC128b<2>.XRES4.B SARP 13.9307f
C267 XA0.CMP_ON a_17462_39772# 0.066018f
C268 XA0.CMP_OP a_2342_40124# 0.066394f
C269 XA6.XA6.Y CK_SAMPLE 0.178114f
C270 XA2.XA8.A VREF 0.028938f
C271 XA6.XA8.A AVDD 1.19556f
C272 XA0.XA1.XA1.MN2.S a_n178_39772# 0.036993f
C273 XA4.XA1.XA1.MP2.S a_11054_40124# 0.04865f
C274 XA2.XA6.Y XA2.DONE 0.014904f
C275 XB2.XA1.Y XB2.M1.G 0.224309f
C276 XA3.CN0 XA6.CN0 0.067216f
C277 XA4.CN0 XA5.CN0 6.498f
C278 XA3.XA1.XA1.MP3.G D<5> 0.014932f
C279 XA2.CN0 XA7.CN0 0.071504f
C280 XA5.XA1.XA1.MP3.S AVDD 0.139093f
C281 XB1.TIE_L XB1.XA2.MP0.G 0.079806f
C282 XA0.CEO a_2342_49100# 0.07472f
C283 XA0.XA11.Y a_974_49100# 0.091063f
C284 a_12422_49452# a_12422_49100# 0.010937f
C285 XDAC1.X16ab.XRES2.B XDAC1.X16ab.XRES1A.B 0.015267f
C286 XA2.XA1.CHL_OP XA0.CMP_OP 0.033149f
C287 XA1.CN1 a_2342_43468# 0.069193f
C288 XA4.EN a_7382_41180# 0.073535f
C289 XA7.CN1 XA8.CN1 0.025286f
C290 XDAC2.XC0.XRES8.B SARN 27.705502f
C291 XA0.CMP_ON XA8.XA1.XA1.MP3.G 0.07295f
C292 XA8.XA10.A XA8.XA6.Y 0.205884f
C293 XA0.XA6.Y XA0.XA8.A 0.527529f
C294 XA5.XA1.XA1.MP3.G a_13574_40476# 0.067588f
C295 XA5.XA1.XA1.MP3.S a_12422_40476# 0.04865f
C296 XA0.XA1.XA1.MP3.S XA0.XA1.XA1.MP2.S 0.050207f
C297 a_3494_46108# CK_SAMPLE 0.07476f
C298 XA7.CN0 SARP 0.036248f
C299 a_2342_46108# D<7> 0.011483f
C300 a_6014_46108# AVDD 0.378183f
C301 XA0.XA1.XA4.MN2.S EN 0.012357f
C302 XA6.XA6.Y XA6.CP0 0.010942f
C303 XA20.XA2.N2 SARP 0.123668f
C304 XA5.CN0 XA0.CMP_OP 0.063388f
C305 XA0.CP0 XA3.CN1 0.147255f
C306 XA1.CP0 XA2.CN1 0.138993f
C307 XA2.CP0 XA1.CN1 0.070579f
C308 XB1.XA3.B m3_7598_1240# 0.024512f
C309 XB1.XA1.MP0.G AVDD 0.518987f
C310 XDAC2.XC128b<2>.XRES16.B XDAC2.XC128b<2>.XRES1A.B 0.467299f
C311 XB2.XA4.GNG m3_16598_4120# 0.0666f
C312 XA0.XA11.Y AVDD 0.712915f
C313 a_22502_48572# XA20.XA10.B 0.034234f
C314 XA3.XA1.XA5.MN2.S XA3.XA1.XA5.MN1.S 0.050207f
C315 XA6.ENO a_18614_39420# 0.082474f
C316 a_16094_41180# a_16094_40828# 0.010937f
C317 XA20.XA1.CK CK_SAMPLE 0.014649f
C318 XA1.ENO VREF 0.879117f
C319 XA0.ENO D<8> 0.101094f
C320 a_974_46988# AVDD 0.395571f
C321 a_9902_39772# a_9902_39420# 0.010937f
C322 XA1.XA1.XA5.MP1.S AVDD 0.102822f
C323 a_16094_42588# EN 0.077363f
C324 XA3.XA6.Y XA3.XA6.MP3.S 0.055045f
C325 a_11054_334# a_11054_n18# 0.010937f
C326 a_7382_46108# XA3.CP0 0.067588f
C327 XA4.CEO XA5.XA10.A 0.019775f
C328 XDAC1.XC128a<1>.XRES1A.B XDAC1.XC32a<0>.XRES1B.B 0.62895f
C329 XA2.XA1.CHL_OP a_4862_41884# 0.040867f
C330 XA1.ENO XA1.XA1.XA1.MN2.S 0.104122f
C331 XA1.CN0 XA1.XA1.XA1.MP3.G 0.013311f
C332 XA4.XA2.A a_11054_42588# 0.129098f
C333 XA0.CMP_ON XA2.XA1.XA5.MN1.S 0.011062f
C334 XA0.CMP_ON a_16094_39772# 0.067588f
C335 XA5.XA1.XA4.MN2.S XA5.XA1.XA4.MN1.S 0.050207f
C336 XA0.CMP_OP a_974_40124# 0.067964f
C337 XA5.XA8.A a_13574_47692# 0.160931f
C338 a_11054_44348# D<4> 0.02026f
C339 a_9614_1918# XB1.M1.G 0.036098f
C340 XA4.CN0 XA4.XA6.MP1.S 0.028026f
C341 XA5.XA1.XA1.MP3.G AVDD 1.05472f
C342 XB1.TIE_L a_9614_2974# 0.03839f
C343 XA0.CEO a_974_49100# 0.015625f
C344 XA4.CEO XA5.XA11.Y 0.293159f
C345 XA0.XA11.Y a_n178_49100# 0.10248f
C346 XA3.CN1 XA0.CMP_ON 0.194649f
C347 XA1.XA1.CHL_OP XA0.CMP_OP 0.03343f
C348 XA6.XA1.CHL_OP XA6.XA2.A 0.133602f
C349 XA0.XA1.CHL_OP a_n178_42588# 0.01727f
C350 XA2.CP0 XA2.XA1.XA4.LCK_N 0.013375f
C351 XDAC1.XC0.XRES4.B SARP 13.930599f
C352 XDAC2.XC32a<0>.XRES2.B SARN 7.01089f
C353 a_17462_48572# AVDD 0.394373f
C354 XA4.XA1.XA4.LCK_N XA4.XA1.XA4.MN1.S 0.030434f
C355 a_11054_48220# XA4.XA6.Y 0.066018f
C356 XA5.XA1.XA1.MP3.G a_12422_40476# 0.096735f
C357 XA0.XA1.XA1.MP3.G XA0.XA1.XA1.MP2.S 0.064105f
C358 XA7.CN0 EN 0.07142f
C359 a_974_46988# XA0.CP1 0.068712f
C360 XA8.XA6.Y a_21134_46108# 0.023316f
C361 XDAC1.XC0.XRES16.B XDAC1.XC64b<1>.XRES16.B 0.010386f
C362 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES8.B 0.029725f
C363 XB1.XA3.B m3_7526_1240# 0.024512f
C364 XB1.XA1.Y AVDD 0.45332f
C365 XA0.CP0 XA2.CN1 0.133733f
C366 a_16094_45228# XA6.XA1.CHL_OP 0.066018f
C367 XA1.CP0 XA1.CN1 0.19197f
C368 XB2.XA4.GNG m3_16526_4120# 0.105547f
C369 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES16.B 0.05157f
C370 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES2.B 0.033713f
C371 XA0.CEO AVDD 1.98375f
C372 a_9902_48572# a_9902_48220# 0.010937f
C373 XA6.ENO a_17462_39420# 0.01235f
C374 XA0.ENO VREF 0.879117f
C375 XA5.ENO D<3> 0.499068f
C376 XA1.XA1.XA4.LCK_N AVDD 0.271288f
C377 a_17462_42588# VREF 0.028416f
C378 XA20.XA4.MP0.S a_22502_45404# 0.023111f
C379 XA1.ENO XA1.XA1.XA1.MP2.S 0.155821f
C380 XA0.ENO XA1.XA1.XA1.MN2.S 0.038148f
C381 XA4.XA2.A a_9902_42588# 0.089492f
C382 XA0.CMP_ON a_14942_39772# 0.066018f
C383 XA0.CMP_OP a_n178_40124# 0.072221f
C384 XA2.XA6.Y VREF 0.078171f
C385 XA4.XA6.Y D<4> 0.039903f
C386 XA6.XA6.Y AVDD 0.864413f
C387 XA4.XA1.XA1.MP3.G a_11054_39420# 0.03422f
C388 XA4.XA1.XA1.MN2.S a_9902_40124# 0.056787f
C389 a_17462_44348# AVDD 0.377363f
C390 a_2342_44348# VREF 0.059568f
C391 a_974_44348# D<8> 0.066018f
C392 XA20.XA2.N1 SARP 0.435464f
C393 XA5.XA8.A a_12422_47692# 0.133834f
C394 XA5.XA6.Y a_13574_47692# 0.017683f
C395 XB2.XA1.Y a_13862_1918# 0.091934f
C396 a_8462_1918# XB1.M1.G 0.072612f
C397 XA8.ENO XA8.CP0 0.08098f
C398 XA4.XA1.XA1.MP3.S AVDD 0.139596f
C399 XA4.CEO XA5.CEO 0.432008f
C400 a_11054_49452# a_11054_49100# 0.010937f
C401 XDAC2.X16ab.XRES2.B XDAC2.X16ab.XRES16.B 0.470901f
C402 XDAC2.X16ab.XRES8.B XDAC2.X16ab.XRES1A.B 0.029729f
C403 XA2.CN1 XA0.CMP_ON 0.192198f
C404 XA0.XA1.CHL_OP XA0.CMP_OP 0.033149f
C405 XA2.ENO a_6014_41180# 0.072087f
C406 XDAC1.XC32a<0>.XRES8.B SARP 27.705599f
C407 a_16094_48572# AVDD 0.394716f
C408 XA0.CMP_OP a_4862_40828# 0.014592f
C409 XA0.CMP_ON XA7.XA1.XA1.MP3.G 0.073013f
C410 XA7.XA10.A XA7.XA9.MN1.S 0.073313f
C411 a_9902_48220# XA4.XA6.Y 0.072725f
C412 XA0.XA1.XA1.MP3.G XA0.XA1.XA1.MN2.S 0.078539f
C413 XA7.XA6.MP1.S D<1> 0.016737f
C414 XA7.CN0 D<8> 0.172519f
C415 a_21134_41884# EN 0.141376f
C416 XA2.XA1.XA4.MP1.S AVDD 0.105303f
C417 XA0.CP0 XA1.CN1 0.137819f
C418 XB1.XA3.B m3_974_2040# 0.0666f
C419 a_14942_45228# XA6.XA1.CHL_OP 0.06825f
C420 XDAC1.XC128b<2>.XRES16.B XDAC1.XC128b<2>.XRES1A.B 0.467299f
C421 a_21134_48572# XA8.XA10.A 0.066018f
C422 a_21134_49452# AVDD 0.46908f
C423 XA3.XA1.XA5.MN2.S XA3.XA1.XA4.LCK_N 0.010898f
C424 XA6.ENO a_16094_39420# 0.010025f
C425 a_14942_41180# a_14942_40828# 0.010937f
C426 XA4.ENO D<3> 0.070845f
C427 a_22502_47164# CK_SAMPLE 0.012715f
C428 XA20.XA1.CK AVDD 3.92726f
C429 a_8534_39772# a_8534_39420# 0.010937f
C430 XA7.XA6.Y a_18614_46988# 0.047651f
C431 a_16094_42588# VREF 0.028416f
C432 a_9614_334# a_9614_n18# 0.010937f
C433 a_6014_46108# XA2.CP0 0.066018f
C434 a_7382_39772# AVDD 0.382762f
C435 XA8.XA1.CHL_OP XA8.XA1.XA5.MN1.S 0.011494f
C436 XA1.XA1.CHL_OP a_3494_41884# 0.040867f
C437 XA7.ENO a_17462_40476# 0.016912f
C438 XDAC2.XC128b<2>.XRES4.B SARN 13.9307f
C439 XA0.CMP_ON a_13574_39772# 0.067588f
C440 XA5.XA6.Y CK_SAMPLE 0.17922f
C441 XA4.XA1.XA1.MP3.G a_9902_39420# 0.023111f
C442 a_21134_40476# a_21134_40124# 0.010937f
C443 a_16094_44348# AVDD 0.377363f
C444 a_974_44348# VREF 0.059568f
C445 XA1.XA8.A XA1.DONE 0.1303f
C446 a_n178_44348# D<8> 0.069545f
C447 XB2.XA1.MP0.G XB2.M1.G 0.036274f
C448 XA2.CN0 XA6.CN0 0.091206f
C449 XA4.XA1.XA1.MP3.G AVDD 1.07016f
C450 XA2.XA1.XA1.MP3.G D<6> 0.017273f
C451 XA4.CEO XA4.XA11.Y 0.158152f
C452 XA1.CN1 XA0.CMP_ON 0.191369f
C453 XA5.XA1.CHL_OP XA5.XA2.A 0.133602f
C454 XA20.XA2.VMR XA0.CMP_OP 0.674482f
C455 XA2.ENO a_4862_41180# 0.068502f
C456 XA0.XA1.XA4.LCK_N a_974_41180# 0.023475f
C457 XA8.XA1.XA4.LCK_N a_19982_41884# 0.031412f
C458 XA0.CMP_OP a_3494_40828# 0.014652f
C459 XA7.XA10.A XA7.XA8.A 0.062692f
C460 XA4.XA1.XA1.MP3.S a_11054_40476# 0.04865f
C461 XA7.CN0 VREF 0.49936f
C462 a_2342_46108# AVDD 0.378183f
C463 a_n178_46108# CK_SAMPLE 0.073189f
C464 XA6.CN0 SARP 0.032152f
C465 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES4.B 0.430615f
C466 XB1.XA3.B m3_830_2040# 0.172147f
C467 XA0.CN0 XA0.XA1.XA4.LCK_N 0.012683f
C468 a_8462_2270# AVDD 0.469157f
C469 XA4.CN0 XA0.CMP_OP 0.06443f
C470 XA20.XA2.CO XA20.XA2.VMR 1.43914f
C471 XA6.ENO XA6.XA1.XA4.LCK_N 0.152052f
C472 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES16.B 0.05157f
C473 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES2.B 0.033713f
C474 a_19982_48572# XA8.XA10.A 0.068275f
C475 a_8534_48572# a_8534_48220# 0.010937f
C476 XA7.CEO XA7.XA6.Y 0.021942f
C477 XA8.ENO CK_SAMPLE 0.130358f
C478 XA4.ENO D<4> 0.431648f
C479 XA7.XA6.Y a_17462_46988# 0.023982f
C480 a_12422_42588# EN 0.078934f
C481 a_4862_46108# XA2.CP0 0.067789f
C482 a_6014_39772# AVDD 0.382569f
C483 XA3.XA11.MP1.S XA3.XA10.Y 0.010335f
C484 XA1.XA1.CHL_OP a_2342_41884# 0.023777f
C485 XDAC1.XC128b<2>.XRES1B.B SARP 3.63755f
C486 XA0.ENO XA0.XA1.XA1.MP2.S 0.150467f
C487 XA3.XA2.A a_8534_42588# 0.091063f
C488 XA0.CMP_ON XA2.XA1.XA4.LCK_N 0.276413f
C489 XA0.CMP_ON a_12422_39772# 0.066018f
C490 XA0.CMP_OP XA8.XA1.XA1.MN2.S 0.024943f
C491 XA5.XA8.A AVDD 1.19556f
C492 XA1.XA8.A VREF 0.028938f
C493 XA8.XA1.XA1.MP3.G a_21134_39772# 0.033843f
C494 XA3.XA1.XA1.MN2.S a_8534_40124# 0.056787f
C495 XA1.XA6.Y XA1.DONE 0.014904f
C496 XA8.XA9.MN1.S XA8.XA8.A 0.010335f
C497 XA20.XA10.A XA20.XA11.MP1.S 0.054658f
C498 XB1.XA1.MP0.G XB1.CKN 0.015687f
C499 XB2.XA1.MP0.G a_15014_1918# 0.067588f
C500 XB1.XA1.Y XB1.XA4.MN1.S 0.011382f
C501 XA7.ENO XA7.CP0 0.08098f
C502 XA3.XA1.XA1.MP3.S AVDD 0.139093f
C503 a_21134_49452# XA8.XA11.Y 0.066018f
C504 a_9902_49452# a_9902_49100# 0.010937f
C505 XDAC1.X16ab.XRES2.B XDAC1.X16ab.XRES16.B 0.470901f
C506 XDAC1.X16ab.XRES8.B XDAC1.X16ab.XRES1A.B 0.029729f
C507 XA20.XA2.CO XA0.CMP_OP 0.144663f
C508 XA20.XA2.VMR a_23654_43116# 0.066661f
C509 XDAC2.XC0.XRES4.B SARN 13.930901f
C510 a_13862_n18# CK_SAMPLE_BSSW 0.011707f
C511 XA7.CN0 XA7.XA1.XA4.LCK_N 0.01537f
C512 XA5.CN1 XA6.CN1 0.025286f
C513 XDAC2.XC1.XRES16.B XDAC2.XC1.XRES1A.B 0.467299f
C514 XA0.XA1.XA4.LCK_N a_n178_41180# 0.060353f
C515 XA0.CMP_ON XA6.XA1.XA1.MP3.G 0.073013f
C516 XA7.XA10.A XA7.XA6.Y 0.205884f
C517 XA4.XA1.XA1.MP3.G a_11054_40476# 0.098305f
C518 XA6.CN0 EN 0.071885f
C519 a_974_46108# AVDD 0.378183f
C520 XA7.CN0 SARN 0.05312f
C521 XA8.XA6.MP3.S D<0> 0.028396f
C522 XA1.ENO XA1.CN0 0.158125f
C523 XA5.XA6.Y XA5.CP0 0.010942f
C524 XA3.XA1.XA4.MP2.S AVDD 0.035519f
C525 XB1.XA3.B m3_7598_2200# 0.024512f
C526 a_13574_45228# XA5.XA1.CHL_OP 0.066679f
C527 XDAC2.XC128b<2>.XRES2.B XDAC2.XC128b<2>.XRES1A.B 0.015267f
C528 XA5.ENO XA6.XA1.XA4.LCK_N 0.339883f
C529 XA3.XA1.XA5.MP2.S XA3.XA1.XA5.MP1.S 0.050207f
C530 XA5.ENO a_14942_39420# 0.071936f
C531 a_13574_41180# a_13574_40828# 0.010937f
C532 XA7.ENO CK_SAMPLE 0.111217f
C533 XA8.ENO DONE 0.041026f
C534 a_22502_47164# AVDD 0.395794f
C535 a_7382_39772# a_7382_39420# 0.010937f
C536 XA0.XA1.XA5.MP1.S AVDD 0.102822f
C537 XA1.XA6.Y XA1.XA6.MN1.S 0.026506f
C538 XA2.XA6.Y XA2.XA6.MP3.S 0.055045f
C539 a_11054_42588# EN 0.077363f
C540 a_8462_334# a_8462_n18# 0.010937f
C541 XA4.CEIN XA3.XA10.A 0.010854f
C542 XA8.XA1.CHL_OP XA8.XA1.XA4.LCK_N 0.204048f
C543 XA0.ENO XA0.XA1.XA1.MN2.S 0.040976f
C544 XA6.ENO a_16094_40476# 0.017441f
C545 XA3.CN1 XA3.XA1.XA4.LCK_N 0.035711f
C546 XA3.XA2.A a_7382_42588# 0.127528f
C547 XA0.CMP_ON XA1.XA1.XA5.MN1.S 0.011178f
C548 XA5.XA1.XA4.MP2.S XA5.XA1.XA4.MP1.S 0.050207f
C549 XA0.CMP_ON a_11054_39772# 0.067588f
C550 XA0.CP1 XDAC1.XC0.XRES16.B 0.031495f
C551 XA0.CMP_OP XA7.XA1.XA1.MN2.S 0.024423f
C552 XA5.XA6.Y AVDD 0.864413f
C553 XA1.XA6.Y VREF 0.078171f
C554 a_19982_40476# a_19982_40124# 0.010937f
C555 XA8.XA1.CHL_OP EN 0.109026f
C556 a_7382_44348# D<5> 0.02026f
C557 XA4.XA8.A a_11054_47692# 0.133834f
C558 XB2.XA1.MP0.G a_13862_1918# 0.071837f
C559 XB1.XA1.MP0.G XB1.XA4.GNG 0.018609f
C560 a_15014_2270# a_15014_1918# 0.010937f
C561 XB1.XA1.Y XB1.CKN 0.200119f
C562 XA0.CP1 a_974_46108# 0.011483f
C563 XA3.XA1.XA1.MP3.G AVDD 1.05472f
C564 XA4.CEIN XA4.XA11.Y 0.220689f
C565 a_21134_49452# XA8.CEO 0.043351f
C566 a_19982_49452# XA8.XA11.Y 0.070936f
C567 XA1.ENO a_3494_41180# 0.06753f
C568 XA4.XA1.CHL_OP XA4.XA2.A 0.133602f
C569 XA20.XA2.CO a_23654_43116# 0.067834f
C570 XA20.XA2.VMR a_22502_43116# 0.078616f
C571 XDAC1.XC0.XRES1B.B SARP 3.64058f
C572 XA1.CP0 XA1.XA1.XA4.LCK_N 0.013291f
C573 XDAC1.XC32a<0>.XRES16.B D<6> 0.018765f
C574 XDAC2.XC32a<0>.XRES8.B SARN 27.705599f
C575 a_12422_48572# AVDD 0.394373f
C576 XA4.XA1.XA1.MP3.G a_9902_40476# 0.066018f
C577 XA6.CN0 D<8> 0.073351f
C578 a_17462_41884# EN 0.143959f
C579 XA0.ENO XA1.CN0 0.058697f
C580 XA2.XA1.XA4.MP2.S AVDD 0.035519f
C581 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES4.B 0.430615f
C582 XB1.XA3.B m3_7526_2200# 0.024512f
C583 a_12422_45228# XA5.XA1.CHL_OP 0.067588f
C584 a_18614_48572# XA7.XA10.A 0.066704f
C585 a_7382_48572# a_7382_48220# 0.010937f
C586 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES8.B 0.477132f
C587 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES2.B 0.015267f
C588 a_17462_49452# AVDD 0.468932f
C589 XA6.ENO CK_SAMPLE 0.111173f
C590 XA8.ENO AVDD 4.23774f
C591 XA4.EN D<5> 0.486956f
C592 XA1.XA6.Y XA1.XA6.MP1.S 0.055045f
C593 a_12422_42588# VREF 0.028416f
C594 XA3.CN0 XA3.XA1.CHL_OP 0.036494f
C595 a_3494_46108# XA1.CP0 0.066219f
C596 XA8.CN0 XA8.CP0 0.676717f
C597 XA0.XA1.CHL_OP a_974_41884# 0.023777f
C598 XA0.CN0 XA0.XA1.XA1.MP3.G 0.017163f
C599 XA0.CMP_ON a_9902_39772# 0.066018f
C600 XA4.XA8.A AVDD 1.19556f
C601 XA4.XA6.Y CK_SAMPLE 0.178114f
C602 XA3.XA6.Y D<5> 0.039903f
C603 XA0.XA8.A VREF 0.028938f
C604 XA3.XA1.XA1.MP3.G a_8534_39420# 0.023111f
C605 XA3.XA1.XA1.MP2.S a_7382_40124# 0.04865f
C606 XA0.XA8.A XA0.DONE 0.1303f
C607 XA8.XA6.Y XA8.XA8.A 0.527529f
C608 XA4.XA8.A a_9902_47692# 0.160931f
C609 XA7.XA1.CHL_OP EN 0.11263f
C610 a_12422_44348# AVDD 0.377363f
C611 XA20.XA2.N1 SARN 0.390202f
C612 XA2.XA1.XA1.MP3.S AVDD 0.139596f
C613 XA6.ENO XA6.CP0 0.08098f
C614 XA1.XA1.XA1.MP3.G D<7> 0.014932f
C615 XA4.CEIN XA4.CEO 0.033943f
C616 a_19982_49452# XA8.CEO 0.023111f
C617 a_8534_49452# a_8534_49100# 0.010937f
C618 XDAC2.X16ab.XRES8.B XDAC2.X16ab.XRES16.B 0.1057f
C619 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES1A.B 0.022835f
C620 XA1.ENO a_2342_41180# 0.073535f
C621 XA20.XA2.CO a_22502_43116# 0.098944f
C622 XDAC1.XC32a<0>.XRES4.B SARP 13.9307f
C623 XDAC1.XC1.XRES16.B XDAC1.XC1.XRES1A.B 0.467299f
C624 a_11054_48572# AVDD 0.394716f
C625 XA0.CMP_OP a_n178_40828# 0.014592f
C626 XA0.CMP_ON XA5.XA1.XA1.MP3.G 0.073013f
C627 XA4.XA1.XA4.LCK_N XA4.XA1.XA4.MN2.S 0.030434f
C628 a_8534_48220# XA3.XA6.Y 0.071154f
C629 XA6.XA10.A XA6.XA8.A 0.062692f
C630 XA8.XA1.XA1.MP3.G XA8.XA1.XA1.MP3.S 0.073693f
C631 XA20.XA4.MP0.S AVDD 0.404908f
C632 XA7.CN0 D<1> 3.2381f
C633 XA6.CN0 VREF 0.496795f
C634 XA8.XA6.MN1.S CK_SAMPLE 0.033706f
C635 a_16094_41884# EN 0.143959f
C636 XB1.XA3.B m3_974_3000# 0.0666f
C637 a_15014_2622# AVDD 0.489453f
C638 XA5.CN0 XA5.XA2.A 0.035115f
C639 XDAC1.XC128b<2>.XRES2.B XDAC1.XC128b<2>.XRES1A.B 0.015267f
C640 a_17462_48572# XA7.XA10.A 0.067588f
C641 a_16094_49452# AVDD 0.468559f
C642 XA4.ENO a_13574_39420# 0.082474f
C643 XA3.CP0 XA3.XA1.XA1.MP3.G 0.016439f
C644 a_12422_41180# a_12422_40828# 0.010937f
C645 XA5.ENO CK_SAMPLE 0.111217f
C646 XA7.ENO AVDD 3.97652f
C647 XA2.ENO D<5> 0.063821f
C648 a_6014_39772# a_6014_39420# 0.010937f
C649 a_21134_47692# a_21134_47340# 0.010937f
C650 XA1.XA1.XA5.MP2.S AVDD 0.038567f
C651 a_11054_42588# VREF 0.028416f
C652 a_15014_686# a_15014_334# 0.010937f
C653 a_2342_46108# XA1.CP0 0.067588f
C654 a_2342_39772# AVDD 0.382762f
C655 XA2.CEO XA3.XA10.A 0.019775f
C656 XDAC2.XC128a<1>.XRES16.B XDAC2.XC128a<1>.XRES1A.B 0.467299f
C657 XA7.XA1.CHL_OP XA7.XA1.XA5.MN1.S 0.011494f
C658 XA0.XA1.CHL_OP a_n178_41884# 0.040867f
C659 XDAC2.XC128b<2>.XRES1B.B SARN 3.63755f
C660 XA2.XA2.A a_6014_42588# 0.129098f
C661 XA0.CMP_ON XA1.XA1.XA4.LCK_N 0.284482f
C662 XA0.CMP_ON a_8534_39772# 0.067588f
C663 XA3.XA1.XA1.MP3.G a_7382_39420# 0.03422f
C664 a_18614_40476# a_18614_40124# 0.010937f
C665 XA8.XA6.Y XA8.XA9.MN1.S 0.023798f
C666 XA6.XA1.CHL_OP EN 0.112859f
C667 a_6014_44348# D<6> 0.02026f
C668 a_11054_44348# AVDD 0.377363f
C669 XA8.XA1.CHL_OP VREF 0.285126f
C670 XA20.XA3.N2 SARN 0.144871f
C671 a_13862_2270# a_13862_1918# 0.010937f
C672 XA2.XA1.XA1.MP3.G AVDD 1.07016f
C673 XA3.CN0 XA5.CN0 0.108912f
C674 XA1.CN0 XA7.CN0 0.158963f
C675 XA4.CEIN XA3.XA11.Y 0.377598f
C676 XA8.XA1.CHL_OP a_19982_43468# 0.010411f
C677 XA3.XA1.CHL_OP XA3.XA2.A 0.133602f
C678 XDAC1.XC0.XRES1B.B D<8> 0.012853f
C679 a_9614_n18# CK_SAMPLE_BSSW 0.011707f
C680 a_21134_44348# XA8.CN1 0.066018f
C681 XA8.XA10.Y VREF 0.014206f
C682 XA7.XA1.XA4.LCK_N a_18614_41884# 0.031412f
C683 XA3.XA1.XA4.LCK_N XA3.XA1.XA4.MN1.S 0.030434f
C684 a_7382_48220# XA3.XA6.Y 0.067588f
C685 XA6.XA10.A XA6.XA9.MN1.S 0.073313f
C686 a_21134_40828# a_21134_40476# 0.010937f
C687 XA0.CP0 XDAC1.XC128b<2>.XRES16.B 0.028741f
C688 XA8.XA6.MP1.S AVDD 0.102754f
C689 XA6.CN0 SARN 0.049024f
C690 XA8.CN0 CK_SAMPLE 0.023396f
C691 XA7.CN0 D<2> 0.142721f
C692 XA8.ENO a_21134_46988# 0.077282f
C693 XA7.XA6.Y a_17462_46108# 0.023316f
C694 XA1.XA1.XA4.MP1.S AVDD 0.105303f
C695 a_11054_45228# XA4.XA1.CHL_OP 0.066018f
C696 XB1.XA3.B m3_830_3000# 0.172147f
C697 XA5.ENO XA5.XA1.XA4.LCK_N 0.154232f
C698 a_6014_48572# a_6014_48220# 0.010937f
C699 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES8.B 0.477132f
C700 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES2.B 0.015267f
C701 XA4.ENO a_12422_39420# 0.01235f
C702 XA4.ENO CK_SAMPLE 0.111173f
C703 XA2.ENO D<6> 0.427123f
C704 XA6.ENO AVDD 4.67622f
C705 XA6.XA6.Y a_16094_46988# 0.023982f
C706 XA0.XA1.XA5.MP2.S AVDD 0.038567f
C707 a_7382_42588# EN 0.078934f
C708 a_974_39772# AVDD 0.382569f
C709 XA2.XA10.Y XA2.XA11.MP1.S 0.010335f
C710 XDAC1.X16ab.XRES1A.B SARP 3.63804f
C711 XA2.XA2.A a_4862_42588# 0.089492f
C712 XA0.CMP_ON a_7382_39772# 0.066018f
C713 XA0.CMP_OP XA6.XA1.XA1.MN2.S 0.024478f
C714 XA4.XA6.Y AVDD 0.864413f
C715 XA2.XA1.XA1.MP2.S a_6014_40124# 0.04865f
C716 XA4.XA6.Y a_9902_47692# 0.017683f
C717 XA5.XA1.CHL_OP EN 0.11263f
C718 XA7.XA1.CHL_OP VREF 0.288305f
C719 XA5.ENO XA5.CP0 0.08098f
C720 XA20.XA1.CKN XA20.XA2.VMR 0.137745f
C721 XA1.XA1.XA1.MP3.S AVDD 0.139093f
C722 a_18614_49452# XA7.XA11.Y 0.069366f
C723 a_7382_49452# a_7382_49100# 0.010937f
C724 XDAC1.X16ab.XRES8.B XDAC1.X16ab.XRES16.B 0.1057f
C725 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES1A.B 0.022835f
C726 XA7.ENO XA8.XA1.XA4.MN2.S 0.012065f
C727 XA0.ENO a_974_41180# 0.072087f
C728 XDAC2.XC0.XRES1B.B SARN 3.65882f
C729 a_19982_44348# XA8.CN1 0.069545f
C730 XA3.CN1 XA4.CN1 0.025642f
C731 XA7.XA10.Y VREF 0.01109f
C732 XDAC2.XC1.XRES2.B XDAC2.XC1.XRES1A.B 0.015267f
C733 XA0.CMP_OP a_19982_41180# 0.086332f
C734 XA0.CMP_ON XA4.XA1.XA1.MP3.G 0.073013f
C735 XA6.XA10.A XA6.XA6.Y 0.205884f
C736 XA3.XA1.XA1.MP3.S a_7382_40476# 0.04865f
C737 XA3.XA1.XA1.MP3.G a_8534_40476# 0.067588f
C738 XA7.XA6.MN1.S CK_SAMPLE 0.053284f
C739 XA7.CN0 D<3> 0.155005f
C740 XA6.XA6.MP1.S D<2> 0.016737f
C741 XA0.ENO XA0.CN0 0.093196f
C742 XA8.ENO a_19982_46988# 0.066245f
C743 XA4.XA6.Y XA4.CP0 0.010942f
C744 a_9902_45228# XA4.XA1.CHL_OP 0.06825f
C745 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128b<2>.XRES1A.B 0.029729f
C746 XA4.ENO XA5.XA1.XA4.LCK_N 0.3401f
C747 XA5.ENO XA6.XA1.XA5.MN2.S 0.010423f
C748 XB1.XA3.B m3_7598_3160# 0.024512f
C749 a_16094_48572# XA6.XA10.A 0.066018f
C750 XA4.ENO a_11054_39420# 0.010025f
C751 a_11054_41180# a_11054_40828# 0.010937f
C752 XA4.EN CK_SAMPLE 0.111217f
C753 XA5.ENO AVDD 3.97532f
C754 a_4862_39772# a_4862_39420# 0.010937f
C755 a_19982_47692# a_19982_47340# 0.010937f
C756 XA6.XA6.Y a_14942_46988# 0.047651f
C757 XA1.XA6.Y XA1.CN0 0.093605f
C758 XA0.XA1.XA4.LCK_N AVDD 0.27148f
C759 a_6014_42588# EN 0.077363f
C760 XB2.XA3.B a_15014_n18# 0.01534f
C761 a_13862_686# a_13862_334# 0.010937f
C762 a_974_46108# XA0.CP0 0.066018f
C763 XA20.XA1.CK a_23654_43996# 0.073227f
C764 XA20.XA1.CKN XA0.CMP_OP 0.01106f
C765 XDAC1.XC128a<1>.XRES16.B XDAC1.XC128a<1>.XRES1A.B 0.467299f
C766 XA8.XA1.CHL_OP XA8.XA1.XA5.MN2.S 0.013533f
C767 XA20.XA2.VMR a_23654_42236# 0.134249f
C768 XA7.XA1.CHL_OP XA7.XA1.XA4.LCK_N 0.204048f
C769 XA5.ENO a_12422_40476# 0.016912f
C770 XA4.XA1.XA4.MP2.S XA4.XA1.XA4.MP1.S 0.050207f
C771 XA0.CMP_ON a_6014_39772# 0.067588f
C772 XA0.CMP_OP XA5.XA1.XA1.MN2.S 0.024423f
C773 XA3.XA6.Y CK_SAMPLE 0.17922f
C774 XA7.XA1.XA1.MP3.G a_17462_39772# 0.033843f
C775 a_17462_40476# a_17462_40124# 0.010937f
C776 XA8.XA1.CHL_OP D<0> 0.193133f
C777 XA4.XA1.CHL_OP EN 0.112859f
C778 XA6.XA1.CHL_OP VREF 0.288305f
C779 XB1.XA1.MP0.G XB1.M1.G 0.036274f
C780 XB2.XA1.MP0.G XB2.XA1.Y 0.22339f
C781 XA20.XA1.CKN XA20.XA2.CO 0.136678f
C782 XA1.XA1.XA1.MP3.G AVDD 1.05472f
C783 XA2.CEO XA3.XA11.Y 0.293159f
C784 a_18614_49452# XA7.CEO 0.024074f
C785 a_17462_49452# XA7.XA11.Y 0.067588f
C786 XA0.ENO a_n178_41180# 0.068502f
C787 XA7.XA1.CHL_OP a_18614_43468# 0.010411f
C788 XA2.XA1.CHL_OP XA2.XA2.A 0.133602f
C789 a_11054_n18# SARP 0.023666f
C790 a_15014_334# CK_SAMPLE_BSSW 0.068023f
C791 a_7382_48572# AVDD 0.394373f
C792 XDAC2.XC32a<0>.XRES4.B SARN 13.9307f
C793 XA0.CMP_OP a_18614_41180# 0.086948f
C794 XA3.XA1.XA1.MP3.G a_7382_40476# 0.096735f
C795 a_19982_40828# a_19982_40476# 0.010937f
C796 XA8.CN0 AVDD 1.33209f
C797 XA6.CN0 D<1> 0.073349f
C798 XA7.XA6.MP1.S CK_SAMPLE 0.022628f
C799 a_12422_41884# EN 0.143959f
C800 a_8462_2622# AVDD 0.491023f
C801 XB1.XA4.GNG m3_974_120# 0.024512f
C802 XA0.CP1 XA0.XA1.XA4.LCK_N 0.015734f
C803 XB1.XA3.B m3_7526_3160# 0.024512f
C804 a_14942_48572# XA6.XA10.A 0.068275f
C805 a_4862_48572# a_4862_48220# 0.010937f
C806 XDAC2.XC32a<0>.XRES16.B XDAC2.XC64a<0>.XRES16.B 0.010386f
C807 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES8.B 0.029725f
C808 a_12422_49452# AVDD 0.468932f
C809 XA2.XA1.XA5.MP2.S XA2.XA1.XA5.MP1.S 0.050207f
C810 XA2.CP0 XA2.XA1.XA1.MP3.G 0.019683f
C811 XA2.ENO CK_SAMPLE 0.111173f
C812 XA1.ENO D<7> 0.486956f
C813 XA4.ENO AVDD 4.67622f
C814 XA2.XA6.Y XA2.XA6.MN3.S 0.089305f
C815 a_7382_42588# VREF 0.028416f
C816 a_n178_46108# XA0.CP0 0.067789f
C817 XA20.XA1.CK a_22502_43996# 0.066018f
C818 XA2.CN0 XA2.XA1.CHL_OP 0.036653f
C819 a_21134_40124# AVDD 0.359431f
C820 XA20.XA2.CO a_23654_42236# 0.023357f
C821 XA20.XA2.VMR a_22502_42236# 0.151031f
C822 XA1.XA2.A a_3494_42588# 0.091063f
C823 XA0.CMP_ON a_4862_39772# 0.066018f
C824 XA2.XA6.Y D<6> 0.039903f
C825 XA3.XA8.A AVDD 1.19556f
C826 XA2.XA1.XA1.MN2.S a_4862_40124# 0.056787f
C827 XA2.XA1.XA1.MP3.G a_6014_39420# 0.03422f
C828 XA3.XA1.CHL_OP EN 0.11263f
C829 a_7382_44348# AVDD 0.377363f
C830 XA5.XA1.CHL_OP VREF 0.288305f
C831 XB1.XA1.Y XB1.M1.G 0.224309f
C832 XB1.XA1.MP0.G a_9614_1918# 0.073407f
C833 a_15014_2270# XB2.XA1.Y 0.030771f
C834 XA1.CN0 XA6.CN0 0.173007f
C835 XA4.ENO XA4.CP0 0.08098f
C836 XA0.CN0 XA7.CN0 0.177906f
C837 XA3.CN0 XA4.CN0 4.14292f
C838 XA2.CN0 XA5.CN0 0.068733f
C839 XA0.XA1.XA1.MP3.S AVDD 0.139596f
C840 a_6014_49452# a_6014_49100# 0.010937f
C841 a_17462_49452# XA7.CEO 0.029627f
C842 XA2.CEO XA4.CEIN 0.432008f
C843 XDAC2.X16ab.XRES8.B XDAC2.X16ab.XRES2.B 0.446669f
C844 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES16.B 0.063821f
C845 XA6.ENO XA7.XA1.XA4.MN2.S 0.012065f
C846 a_13862_334# CK_SAMPLE_BSSW 0.078536f
C847 a_18614_44348# XA7.CN1 0.067974f
C848 XA2.CN1 XA3.CN1 1.73981f
C849 XDAC1.XC1.XRES2.B XDAC1.XC1.XRES1A.B 0.015267f
C850 a_6014_48572# AVDD 0.394716f
C851 XDAC1.XC32a<0>.XRES1B.B SARP 3.63755f
C852 XA0.CMP_ON XA3.XA1.XA1.MP3.G 0.073013f
C853 XA3.XA1.XA4.LCK_N XA3.XA1.XA4.MN2.S 0.030434f
C854 XA5.XA10.A XA5.XA9.MN1.S 0.073313f
C855 XA7.XA1.XA1.MP3.G XA7.XA1.XA1.MP3.S 0.073693f
C856 XA6.CN0 D<2> 1.94095f
C857 XA5.CN0 SARP 0.032152f
C858 XA7.ENO a_18614_46988# 0.067815f
C859 a_11054_41884# EN 0.143959f
C860 XA0.XA1.XA4.MP1.S AVDD 0.105303f
C861 a_8534_45228# XA3.XA1.CHL_OP 0.066679f
C862 XA4.CN0 XA4.XA2.A 0.035589f
C863 XA3.CN0 XA0.CMP_OP 0.055878f
C864 XA4.ENO XA5.XA1.XA5.MN2.S 0.010423f
C865 XB2.XA2.MP0.G AVDD 0.809596f
C866 XB1.XA4.GNG m3_830_120# 0.049023f
C867 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128b<2>.XRES1A.B 0.029729f
C868 XB1.XA3.B m3_974_3960# 0.0666f
C869 a_11054_49452# AVDD 0.468559f
C870 XA4.EN a_9902_39420# 0.071936f
C871 XA0.CMP_OP a_22502_42236# 0.011396f
C872 XA2.CN0 XDAC2.X16ab.XRES16.B 0.018342f
C873 a_9902_41180# a_9902_40828# 0.010937f
C874 XA1.ENO CK_SAMPLE 0.111217f
C875 XA0.ENO D<7> 0.063821f
C876 XA4.EN AVDD 3.97532f
C877 a_3494_39772# a_3494_39420# 0.010937f
C878 a_18614_47692# a_18614_47340# 0.010937f
C879 a_21134_42588# AVDD 0.376424f
C880 a_6014_42588# VREF 0.028416f
C881 a_12422_686# a_12422_334# 0.010937f
C882 XA8.ENO XA0.CMP_ON 0.297242f
C883 XA1.CEO XA1.XA10.A 0.010854f
C884 XDAC2.XC128a<1>.XRES2.B XDAC2.XC128a<1>.XRES1A.B 0.015267f
C885 XA1.XA2.A a_2342_42588# 0.127528f
C886 XA7.XA1.CHL_OP XA7.XA1.XA5.MN2.S 0.013533f
C887 XA20.XA2.CO a_22502_42236# 0.035145f
C888 XA4.ENO a_11054_40476# 0.017441f
C889 XDAC2.X16ab.XRES1A.B SARN 3.63804f
C890 XA0.CMP_ON XA0.XA1.XA5.MN1.S 0.011062f
C891 XA0.CMP_ON a_3494_39772# 0.067588f
C892 XA3.XA6.Y AVDD 0.864413f
C893 a_16094_40476# a_16094_40124# 0.010937f
C894 XA2.XA1.XA1.MP3.G a_4862_39420# 0.023111f
C895 XA3.XA8.A a_8534_47692# 0.160931f
C896 XA2.XA1.CHL_OP EN 0.112859f
C897 a_2342_44348# D<7> 0.02026f
C898 a_6014_44348# AVDD 0.377363f
C899 XA4.XA1.CHL_OP VREF 0.288305f
C900 XA7.XA1.CHL_OP D<1> 0.209177f
C901 XB1.XA1.Y a_9614_1918# 0.090364f
C902 a_13862_2270# XB2.XA1.Y 0.015779f
C903 XB1.XA1.MP0.G a_8462_1918# 0.066018f
C904 XA0.XA1.XA1.MP3.G AVDD 1.07017f
C905 XA2.CEO XA2.XA11.Y 0.158152f
C906 XA1.XA1.CHL_OP XA1.XA2.A 0.133602f
C907 a_17462_44348# XA7.CN1 0.067588f
C908 XA1.CN1 XA3.CN1 0.216451f
C909 XA6.XA10.Y VREF 0.011196f
C910 XA5.XA10.A XA5.XA8.A 0.062692f
C911 a_6014_48220# XA2.XA6.Y 0.066018f
C912 XA2.XA1.XA1.MP3.S a_6014_40476# 0.04865f
C913 a_18614_40828# a_18614_40476# 0.010937f
C914 XA6.CN0 D<3> 0.152644f
C915 XA7.XA6.MP1.S AVDD 0.092671f
C916 XA5.CN0 EN 0.071169f
C917 a_22502_46812# CK_SAMPLE 0.013762f
C918 a_23654_39420# a_23654_39068# 0.010937f
C919 XA7.ENO a_17462_46988# 0.075712f
C920 XA6.XA6.Y a_16094_46108# 0.023316f
C921 XDAC2.XC0.XRES1A.B XDAC2.XC64b<1>.XRES1B.B 0.62895f
C922 a_7382_45228# XA3.XA1.CHL_OP 0.067588f
C923 XB1.XA4.GNG m3_7598_280# 0.105547f
C924 XB1.XA3.B m3_830_3960# 0.172147f
C925 a_13574_48572# XA5.XA10.A 0.066704f
C926 a_3494_48572# a_3494_48220# 0.010937f
C927 XDAC1.XC32a<0>.XRES16.B XDAC1.XC64a<0>.XRES16.B 0.010386f
C928 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES8.B 0.029725f
C929 XA2.XA1.XA4.LCK_N XA2.XA1.XA5.MN1.S 0.030434f
C930 XA0.ENO CK_SAMPLE 0.111173f
C931 XA2.ENO AVDD 4.67622f
C932 a_2342_42588# EN 0.078934f
C933 XA7.ENO XA0.CMP_ON 1.18395f
C934 XA1.XA11.MP1.S XA1.XA10.Y 0.010335f
C935 XA0.CP1 XA0.XA1.XA1.MP3.G 0.017273f
C936 XDAC1.X16ab.XRES16.B SARP 55.2956f
C937 XA0.CMP_OP XA4.XA1.XA1.MN2.S 0.024478f
C938 XA0.CMP_ON a_2342_39772# 0.066018f
C939 XA2.XA6.Y CK_SAMPLE 0.178114f
C940 XA2.XA8.A AVDD 1.19556f
C941 XA1.XA1.XA1.MN2.S a_3494_40124# 0.056787f
C942 XA6.XA1.XA1.MP3.G a_16094_39772# 0.033843f
C943 XA3.XA8.A a_7382_47692# 0.133834f
C944 XA3.XA6.Y a_8534_47692# 0.017683f
C945 XA7.XA8.A XA7.XA9.MN1.S 0.010335f
C946 XA7.XA6.Y XA8.XA6.Y 0.046858f
C947 XA1.XA1.CHL_OP EN 0.11263f
C948 XA3.XA1.CHL_OP VREF 0.288305f
C949 a_9614_2270# a_9614_1918# 0.010937f
C950 XA4.EN XA3.CP0 0.173089f
C951 a_23654_40828# AVDD 0.024826f
C952 a_4862_49452# a_4862_49100# 0.010937f
C953 a_16094_49452# XA6.XA11.Y 0.066018f
C954 XDAC1.X16ab.XRES8.B XDAC1.X16ab.XRES2.B 0.446669f
C955 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES16.B 0.063821f
C956 XA1.CN1 XA2.CN1 3.3766f
C957 a_12422_334# SAR_IN 0.061868f
C958 a_12422_n18# SARN 0.023465f
C959 XA5.XA10.Y VREF 0.01109f
C960 XDAC2.XC1.XRES2.B XDAC2.XC1.XRES16.B 0.470901f
C961 XDAC2.XC1.XRES8.B XDAC2.XC1.XRES1A.B 0.029729f
C962 XA0.CMP_OP a_14942_41180# 0.085247f
C963 XA0.CMP_ON XA2.XA1.XA1.MP3.G 0.073013f
C964 XA5.XA10.A XA5.XA6.Y 0.205884f
C965 a_4862_48220# XA2.XA6.Y 0.072725f
C966 XA2.XA1.XA1.MP3.G a_6014_40476# 0.098305f
C967 XA5.CN0 D<8> 0.073419f
C968 XA8.XA6.MP3.S CK_SAMPLE 0.016391f
C969 a_23654_46812# AVDD 0.024826f
C970 XA3.XA6.Y XA3.CP0 0.010942f
C971 XA1.XA1.XA4.MP2.S AVDD 0.035519f
C972 XB1.XA4.GNG m3_7526_280# 0.0666f
C973 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES1A.B 0.022835f
C974 XB1.XA3.B m3_7598_4120# 0.024512f
C975 a_12422_48572# XA5.XA10.A 0.067588f
C976 XA2.ENO a_8534_39420# 0.082474f
C977 XA1.CP0 XA1.XA1.XA1.MP3.G 0.016439f
C978 a_8534_41180# a_8534_40828# 0.010937f
C979 XA1.ENO AVDD 3.97532f
C980 a_2342_39772# a_2342_39420# 0.010937f
C981 XA5.XA6.Y a_13574_46988# 0.047651f
C982 a_17462_47692# a_17462_47340# 0.010937f
C983 a_974_42588# EN 0.077363f
C984 a_11054_686# a_11054_334# 0.010937f
C985 XA7.CN0 XA7.CP0 0.796454f
C986 XA6.ENO XA0.CMP_ON 1.03137f
C987 a_17462_40124# AVDD 0.3588f
C988 XA0.CEO XA1.XA10.A 0.019775f
C989 XDAC1.XC128a<1>.XRES2.B XDAC1.XC128a<1>.XRES1A.B 0.015267f
C990 XA0.XA2.A a_974_42588# 0.129098f
C991 XA2.CN1 XA2.XA1.XA4.LCK_N 0.033627f
C992 XDAC1.XC1.XRES1A.B SARP 3.63777f
C993 XA0.CMP_OP XA3.XA1.XA1.MN2.S 0.024423f
C994 XA4.XA1.XA4.MN2.S XA4.XA1.XA4.MN1.S 0.050207f
C995 XA0.CMP_ON a_974_39772# 0.067588f
C996 a_14942_40476# a_14942_40124# 0.010937f
C997 XA7.XA6.Y XA7.XA9.MN1.S 0.023798f
C998 XA6.XA1.CHL_OP D<2> 0.209422f
C999 XA0.XA1.CHL_OP EN 0.242472f
C1000 XA2.XA1.CHL_OP VREF 0.288305f
C1001 XA20.XA2.VMR SARP 0.122801f
C1002 a_15014_2270# XB2.XA1.MP0.G 0.066018f
C1003 XA2.ENO XA3.CP0 0.061526f
C1004 XA2.CN0 XA4.CN0 0.068518f
C1005 XA0.CN0 XA6.CN0 0.188403f
C1006 a_22502_40828# AVDD 0.502735f
C1007 a_14942_49452# XA6.XA11.Y 0.070936f
C1008 a_16094_49452# XA6.CEO 0.040807f
C1009 XA1.CEO XA2.XA11.Y 0.220689f
C1010 XA6.XA1.CHL_OP a_14942_43468# 0.010411f
C1011 XA0.XA1.CHL_OP XA0.XA2.A 0.133602f
C1012 XA0.CP0 XA0.XA1.XA4.LCK_N 0.013375f
C1013 a_16094_44348# XA6.CN1 0.066018f
C1014 a_9614_334# CK_SAMPLE_BSSW 0.080106f
C1015 a_2342_48572# AVDD 0.394373f
C1016 XDAC2.XC32a<0>.XRES1B.B SARN 3.63755f
C1017 XA0.CMP_OP a_13574_41180# 0.086948f
C1018 XA2.XA1.XA1.MP3.G a_4862_40476# 0.066018f
C1019 a_17462_40828# a_17462_40476# 0.010937f
C1020 XA4.CN0 SARP 0.032152f
C1021 XA5.CN0 VREF 0.49936f
C1022 XA7.CN0 CK_SAMPLE 0.075434f
C1023 a_22502_46812# AVDD 0.502744f
C1024 a_22502_39420# a_22502_39068# 0.010937f
C1025 XA6.ENO a_16094_46988# 0.077282f
C1026 a_7382_41884# EN 0.143959f
C1027 XA0.XA1.XA4.MP2.S AVDD 0.035519f
C1028 XDAC1.XC0.XRES1A.B XDAC1.XC64b<1>.XRES1B.B 0.62895f
C1029 a_6014_45228# XA2.XA1.CHL_OP 0.066018f
C1030 XA2.CN0 XA0.CMP_OP 0.057021f
C1031 a_15014_2974# AVDD 0.472782f
C1032 XB1.XA4.GNG m3_974_1080# 0.024512f
C1033 XB1.XA3.B m3_7526_4120# 0.024512f
C1034 a_2342_48572# a_2342_48220# 0.010937f
C1035 a_7382_49452# AVDD 0.468932f
C1036 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES4.B 0.430615f
C1037 XA2.ENO a_7382_39420# 0.01235f
C1038 XA5.CEO XA5.XA6.Y 0.021942f
C1039 XA0.ENO AVDD 4.67625f
C1040 XA5.XA6.Y a_12422_46988# 0.023982f
C1041 XA1.XA6.Y XA1.XA6.MN3.S 0.089305f
C1042 a_n178_42588# EN 0.078848f
C1043 a_17462_42588# AVDD 0.376544f
C1044 a_2342_42588# VREF 0.028416f
C1045 XA8.ENO XA8.CN1 0.083825f
C1046 XA5.ENO XA0.CMP_ON 1.18612f
C1047 a_16094_40124# AVDD 0.358987f
C1048 XA6.XA1.CHL_OP XA6.XA1.XA5.MN1.S 0.011494f
C1049 XA0.CMP_ON XA0.XA1.XA4.LCK_N 0.276252f
C1050 XA0.XA2.A a_n178_42588# 0.089492f
C1051 XA0.CMP_ON a_n178_39772# 0.066018f
C1052 XA2.XA6.Y AVDD 0.864413f
C1053 XA1.XA6.Y D<7> 0.039903f
C1054 XA1.XA1.XA1.MP2.S a_2342_40124# 0.04865f
C1055 XA1.XA1.XA1.MP3.G a_3494_39420# 0.023111f
C1056 XA7.XA6.Y XA7.XA8.A 0.527529f
C1057 a_2342_44348# AVDD 0.377363f
C1058 XA0.XA1.CHL_OP D<8> 0.529833f
C1059 XA1.XA1.CHL_OP VREF 0.288305f
C1060 a_8462_2270# a_8462_1918# 0.010937f
C1061 a_13862_2270# XB2.XA1.MP0.G 0.099734f
C1062 XA2.ENO XA2.CP0 0.111184f
C1063 XA3.CN0 XA3.XA6.MP1.S 0.028026f
C1064 a_21134_40828# AVDD 0.407021f
C1065 a_3494_49452# a_3494_49100# 0.010937f
C1066 a_14942_49452# XA6.CEO 0.023111f
C1067 XA1.CEO XA2.CEO 0.033943f
C1068 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES2.B 0.033713f
C1069 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES16.B 0.05157f
C1070 XA6.CN0 XA6.XA1.XA4.LCK_N 0.015589f
C1071 a_14942_44348# XA6.CN1 0.069545f
C1072 a_11054_334# SAR_IP 0.061868f
C1073 a_8462_334# CK_SAMPLE_BSSW 0.066453f
C1074 a_974_48572# AVDD 0.394716f
C1075 XDAC1.XC1.XRES2.B XDAC1.XC1.XRES16.B 0.470901f
C1076 XDAC1.XC1.XRES8.B XDAC1.XC1.XRES1A.B 0.029729f
C1077 XDAC1.XC128a<1>.XRES1A.B SARP 3.63804f
C1078 XA0.CMP_ON XA1.XA1.XA1.MP3.G 0.073013f
C1079 XA4.XA10.A XA4.XA8.A 0.062692f
C1080 XA6.XA1.XA1.MP3.G XA6.XA1.XA1.MP3.S 0.073693f
C1081 XA5.CN0 SARN 0.049024f
C1082 XA7.XA6.MP3.S D<1> 0.028396f
C1083 XA6.XA6.MP1.S CK_SAMPLE 0.022425f
C1084 XA4.CN0 EN 0.071817f
C1085 XA8.XA6.MP3.S AVDD 0.104402f
C1086 XA6.ENO a_14942_46988# 0.066245f
C1087 XA0.ENO XA0.CP1 0.427123f
C1088 a_6014_41884# EN 0.143959f
C1089 a_4862_45228# XA2.XA1.CHL_OP 0.06825f
C1090 XB1.XA4.GNG m3_830_1080# 0.049023f
C1091 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES1A.B 0.022835f
C1092 a_11054_48572# XA4.XA10.A 0.066018f
C1093 a_6014_49452# AVDD 0.468559f
C1094 XA2.ENO a_6014_39420# 0.010025f
C1095 XA8.ENO a_21134_39772# 0.045171f
C1096 XA0.CMP_OP XA8.XA1.XA4.LCK_N 0.387059f
C1097 a_7382_41180# a_7382_40828# 0.010937f
C1098 a_974_39772# a_974_39420# 0.010937f
C1099 a_16094_47692# a_16094_47340# 0.010937f
C1100 XA20.XA10.A XA20.XA1.CK 0.024853f
C1101 XA1.XA6.Y XA1.XA6.MP3.S 0.055045f
C1102 XA0.CMP_OP EN 1.27092f
C1103 a_974_42588# VREF 0.028416f
C1104 a_16094_42588# AVDD 0.376544f
C1105 XB2.XA3.B a_15014_334# 0.011407f
C1106 a_9614_686# a_9614_334# 0.010937f
C1107 XA8.CN0 a_21134_46108# 0.103403f
C1108 XA4.ENO XA0.CMP_ON 1.03123f
C1109 XDAC2.XC128a<1>.XRES2.B XDAC2.XC128a<1>.XRES16.B 0.470901f
C1110 XDAC2.XC128a<1>.XRES8.B XDAC2.XC128a<1>.XRES1A.B 0.029729f
C1111 XA4.EN a_7382_40476# 0.016912f
C1112 XDAC2.X16ab.XRES16.B SARN 55.2956f
C1113 XA0.CMP_ON a_21134_40124# 0.066018f
C1114 XA1.XA6.Y CK_SAMPLE 0.17922f
C1115 XA0.XA6.Y a_n178_47340# 0.011912f
C1116 a_13574_40476# a_13574_40124# 0.010937f
C1117 XA1.XA1.XA1.MP3.G a_2342_39420# 0.03422f
C1118 XA5.XA1.CHL_OP D<3> 0.209177f
C1119 XA2.XA8.A a_6014_47692# 0.133834f
C1120 a_974_44348# AVDD 0.377363f
C1121 XA0.XA1.CHL_OP VREF 0.288305f
C1122 XA1.CEO XA1.XA11.Y 0.377598f
C1123 XA5.XA1.CHL_OP a_13574_43468# 0.010411f
C1124 a_11054_334# SARP 0.037284f
C1125 a_15014_686# CK_SAMPLE_BSSW 0.066018f
C1126 XA4.XA10.Y VREF 0.011196f
C1127 XA4.XA10.A XA4.XA9.MN1.S 0.073313f
C1128 a_16094_40828# a_16094_40476# 0.010937f
C1129 XA4.CN0 D<8> 0.074539f
C1130 XA5.XA6.MP1.S D<3> 0.016737f
C1131 XA7.CN0 AVDD 4.65707f
C1132 XA6.XA6.MN1.S CK_SAMPLE 0.050648f
C1133 a_21134_39420# a_21134_39068# 0.010937f
C1134 XA20.XA2.N2 AVDD 0.33734f
C1135 XA8.CP0 XA8.XA1.CHL_OP 0.731503f
C1136 XA4.ENO XA4.XA1.XA4.LCK_N 0.152052f
C1137 a_15014_3326# AVDD 0.450704f
C1138 XB1.XA4.GNG m3_7598_1240# 0.105547f
C1139 a_9902_48572# XA4.XA10.A 0.068275f
C1140 a_974_48572# a_974_48220# 0.010937f
C1141 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES4.B 0.430615f
C1142 XA2.XA1.XA5.MN2.S XA2.XA1.XA5.MN1.S 0.050207f
C1143 XA0.CP0 XA0.XA1.XA1.MP3.G 0.019683f
C1144 a_21134_47340# AVDD 0.390024f
C1145 XA8.XA8.A XA8.ENO 0.143506f
C1146 XA0.CMP_OP D<8> 0.223336f
C1147 XA20.XA10.A a_23654_47164# 0.07154f
C1148 XB1.XA3.B a_8462_n18# 0.01534f
C1149 XA7.ENO XA7.CN1 0.083825f
C1150 XA4.EN XA0.CMP_ON 1.18612f
C1151 XA0.CP1 a_974_44348# 0.02026f
C1152 XA0.XA10.Y XA0.XA11.MP1.S 0.010335f
C1153 XDAC1.X16ab.XRES2.B SARP 7.01089f
C1154 XDAC2.XC1.XRES1A.B SARN 3.63777f
C1155 XA0.CMP_OP XA2.XA1.XA1.MN2.S 0.024478f
C1156 XA0.CMP_ON a_19982_40124# 0.074163f
C1157 XA1.XA8.A AVDD 1.19556f
C1158 XA0.XA1.XA1.MP2.S a_974_40124# 0.04865f
C1159 XA2.XA8.A a_4862_47692# 0.160931f
C1160 XA1.ENO XA1.CP0 0.173089f
C1161 a_2342_49452# a_2342_49100# 0.010937f
C1162 a_13574_49452# XA5.XA11.Y 0.069366f
C1163 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES2.B 0.033713f
C1164 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES16.B 0.05157f
C1165 a_13574_44348# XA5.CN1 0.067974f
C1166 a_13862_686# CK_SAMPLE_BSSW 0.072629f
C1167 XA3.XA10.Y VREF 0.01109f
C1168 XDAC2.XC1.XRES8.B XDAC2.XC1.XRES16.B 0.1057f
C1169 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES1A.B 0.022835f
C1170 XA0.CMP_OP a_9902_41180# 0.085247f
C1171 XA0.CMP_ON XA0.XA1.XA1.MP3.G 0.072852f
C1172 XA4.XA10.A XA4.XA6.Y 0.205884f
C1173 a_3494_48220# XA1.XA6.Y 0.071154f
C1174 XA1.XA1.XA1.MP3.S a_2342_40476# 0.04865f
C1175 XA1.XA1.XA1.MP3.G a_3494_40476# 0.067588f
C1176 XA5.CN0 D<1> 0.07328f
C1177 XA4.CN0 VREF 0.496795f
C1178 XA6.XA6.MP3.S D<2> 0.028396f
C1179 XA6.XA6.MP1.S AVDD 0.092671f
C1180 XA6.CN0 CK_SAMPLE 0.075021f
C1181 a_21134_41884# AVDD 0.397696f
C1182 XA2.XA6.Y XA2.CP0 0.010942f
C1183 XA5.ENO a_13574_46988# 0.067815f
C1184 a_3494_45228# XA1.XA1.CHL_OP 0.066679f
C1185 XA4.EN XA4.XA1.XA4.LCK_N 0.339883f
C1186 XB1.XA4.GNG m3_7526_1240# 0.0666f
C1187 XA1.ENO a_4862_39420# 0.071936f
C1188 XA7.ENO a_19982_39772# 0.085451f
C1189 XA8.XA2.A XA8.XA1.XA5.MP2.S 0.050207f
C1190 a_6014_41180# a_6014_40828# 0.010937f
C1191 a_n178_39772# a_n178_39420# 0.010937f
C1192 XA20.XA10.A a_22502_47164# 0.066018f
C1193 a_14942_47692# a_14942_47340# 0.010937f
C1194 a_8462_686# a_8462_334# 0.010937f
C1195 XA7.CN0 XA3.CP0 0.024041f
C1196 XA2.ENO XA0.CMP_ON 1.03123f
C1197 XA6.CN0 XA6.CP0 0.800576f
C1198 a_12422_40124# AVDD 0.3588f
C1199 XB1.TIE_L XA0.XA11.MP1.S 0.010502f
C1200 XDAC1.XC128a<1>.XRES2.B XDAC1.XC128a<1>.XRES16.B 0.470901f
C1201 XDAC1.XC128a<1>.XRES8.B XDAC1.XC128a<1>.XRES1A.B 0.029729f
C1202 XA6.XA1.CHL_OP XA6.XA1.XA4.LCK_N 0.204048f
C1203 XA1.CN1 XA1.XA1.XA4.LCK_N 0.035711f
C1204 XA2.ENO a_6014_40476# 0.017441f
C1205 XA8.ENO XA8.XA1.XA1.MP3.S 0.076247f
C1206 XDAC1.XC1.XRES16.B SARP 55.2953f
C1207 XA0.CMP_OP XA1.XA1.XA1.MN2.S 0.024423f
C1208 XA3.XA1.XA4.MN2.S XA3.XA1.XA4.MN1.S 0.050207f
C1209 XA0.CMP_ON a_18614_40124# 0.072592f
C1210 XA1.XA6.Y AVDD 0.864413f
C1211 a_12422_40476# a_12422_40124# 0.010937f
C1212 XA5.XA1.XA1.MP3.G a_12422_39772# 0.033843f
C1213 XA4.XA1.CHL_OP D<4> 0.209422f
C1214 XA20.XA2.CO VREF 0.030275f
C1215 XA20.XA2.N1 AVDD 0.618791f
C1216 XA20.XA2.VMR SARN 0.052367f
C1217 a_12422_2446# a_12422_2094# 0.010937f
C1218 XA1.CN0 XA5.CN0 0.152661f
C1219 a_17462_40828# AVDD 0.407021f
C1220 XA0.ENO XA1.CP0 0.061526f
C1221 a_12422_49452# XA5.XA11.Y 0.067588f
C1222 a_13574_49452# XA5.CEO 0.024074f
C1223 XA0.CEO XA1.XA11.Y 0.293159f
C1224 a_12422_44348# XA5.CN1 0.067588f
C1225 a_22502_48924# AVDD 0.452052f
C1226 XA0.XA6.Y XA0.XA9.MN1.S 0.023798f
C1227 XDAC2.XC128a<1>.XRES1A.B SARN 3.63804f
C1228 XA6.XA1.XA4.LCK_N a_14942_41884# 0.031412f
C1229 XA0.CMP_OP a_8534_41180# 0.086948f
C1230 a_2342_48220# XA1.XA6.Y 0.067588f
C1231 XA1.XA1.XA1.MP3.G a_2342_40476# 0.096735f
C1232 a_14942_40828# a_14942_40476# 0.010937f
C1233 XA8.XA6.MN3.S CK_SAMPLE 0.044153f
C1234 XA4.CN0 SARN 0.048999f
C1235 XA5.CN0 D<2> 0.066074f
C1236 a_19982_39420# a_19982_39068# 0.010937f
C1237 a_21134_47340# a_21134_46988# 0.010937f
C1238 XA5.ENO a_12422_46988# 0.075712f
C1239 a_2342_41884# EN 0.143959f
C1240 XA5.XA6.Y a_12422_46108# 0.023316f
C1241 a_2342_45228# XA1.XA1.CHL_OP 0.067588f
C1242 XA7.CP0 XA7.XA1.CHL_OP 0.729665f
C1243 XB1.XA2.MP0.G AVDD 0.809596f
C1244 XB1.XA4.GNG m3_974_2040# 0.024512f
C1245 a_8534_48572# XA3.XA10.A 0.066704f
C1246 a_n178_48572# a_n178_48220# 0.010937f
C1247 a_2342_49452# AVDD 0.468932f
C1248 XA0.CMP_OP XA7.XA1.XA4.LCK_N 0.383512f
C1249 XA8.XA1.CHL_OP XA8.XA1.XA4.MP2.S 0.050207f
C1250 XA4.XA6.Y a_11054_46988# 0.023982f
C1251 XA8.XA2.A EN 0.166272f
C1252 a_12422_42588# AVDD 0.376544f
C1253 XA1.CN0 XA1.XA1.CHL_OP 0.036494f
C1254 XA6.ENO XA6.CN1 0.083825f
C1255 XA1.ENO XA0.CMP_ON 1.18612f
C1256 a_11054_40124# AVDD 0.358987f
C1257 XB1.TIE_L XA0.XA10.Y 0.300886f
C1258 XA8.ENO XA8.XA1.XA1.MP3.G 0.328206f
C1259 XA0.CMP_ON a_17462_40124# 0.067588f
C1260 XA8.XA1.XA4.LCK_N a_21134_41180# 0.023475f
C1261 XA0.XA8.A AVDD 1.19559f
C1262 XA0.XA1.XA1.MN2.S a_n178_40124# 0.056787f
C1263 XA0.XA1.XA1.MP3.G a_974_39420# 0.03422f
C1264 a_21134_45228# VREF 0.059517f
C1265 XA2.XA6.Y a_4862_47692# 0.017683f
C1266 XA20.XA3.N2 AVDD 0.32365f
C1267 XA20.XA2.CO SARN 0.202607f
C1268 XA6.XA9.MN1.S XA6.XA8.A 0.010335f
C1269 a_16094_40828# AVDD 0.407021f
C1270 XA0.ENO XA0.CP0 0.111184f
C1271 a_21134_41180# EN 0.074258f
C1272 a_974_49452# a_974_49100# 0.010937f
C1273 a_12422_49452# XA5.CEO 0.029627f
C1274 XA0.CEO XA1.CEO 0.432008f
C1275 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES8.B 0.477132f
C1276 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES2.B 0.015267f
C1277 XA5.ENO XA6.XA1.XA4.MN2.S 0.012065f
C1278 a_12422_334# SARN 0.037174f
C1279 a_12422_686# SAR_IN 0.060109f
C1280 XDAC1.XC1.XRES8.B XDAC1.XC1.XRES16.B 0.1057f
C1281 XA8.XA11.MP1.S AVDD 0.118946f
C1282 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES1A.B 0.022835f
C1283 XB1.TIE_L CK_SAMPLE_BSSW 7.03218f
C1284 XDAC1.XC128a<1>.XRES16.B SARP 55.2956f
C1285 XA3.CN1 XA3.XA1.XA1.MP3.G 0.012023f
C1286 XA3.XA10.A XA3.XA9.MN1.S 0.073313f
C1287 XA5.XA1.XA1.MP3.G XA5.XA1.XA1.MP3.S 0.073693f
C1288 XA7.XA6.MN3.S CK_SAMPLE 0.028234f
C1289 XA6.CN0 AVDD 4.3763f
C1290 XA5.CN0 D<3> 1.85159f
C1291 a_974_41884# EN 0.143959f
C1292 XA3.CN0 XA3.XA2.A 0.02751f
C1293 XB1.XA4.GNG m3_830_2040# 0.049023f
C1294 a_974_49452# AVDD 0.468559f
C1295 a_7382_48572# XA3.XA10.A 0.067588f
C1296 XB1.TIE_L XA0.XA6.Y 0.010239f
C1297 XA0.ENO a_3494_39420# 0.082474f
C1298 XA6.ENO a_18614_39772# 0.082231f
C1299 XA7.ENO a_17462_39772# 0.044989f
C1300 XA1.XA1.XA4.LCK_N XA1.XA1.XA5.MN1.S 0.030434f
C1301 XA2.XA1.XA5.MN2.S XA2.XA1.XA4.LCK_N 0.010898f
C1302 SAR_IN CK_SAMPLE_BSSW 0.016648f
C1303 a_4862_41180# a_4862_40828# 0.010937f
C1304 XA20.XA1.CKN SARP 0.45433f
C1305 a_17462_47340# AVDD 0.390024f
C1306 a_21134_40124# a_21134_39772# 0.010937f
C1307 XA4.XA6.Y a_9902_46988# 0.047651f
C1308 XA8.XA6.Y XA8.ENO 0.051206f
C1309 a_13574_47692# a_13574_47340# 0.010937f
C1310 XA7.XA2.A EN 0.166192f
C1311 a_11054_42588# AVDD 0.376544f
C1312 XA0.ENO XA0.CMP_ON 1.03107f
C1313 XDAC2.XC128a<1>.XRES8.B XDAC2.XC128a<1>.XRES16.B 0.1057f
C1314 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES1A.B 0.022835f
C1315 XA5.XA1.CHL_OP XA5.XA1.XA5.MN1.S 0.011494f
C1316 a_21134_43468# XA8.XA2.A 0.066256f
C1317 XA7.ENO XA8.XA1.XA1.MP3.G 0.031869f
C1318 XDAC2.X16ab.XRES2.B SARN 7.01089f
C1319 XA0.CMP_ON a_16094_40124# 0.066018f
C1320 XA8.XA1.XA4.LCK_N a_19982_41180# 0.060353f
C1321 a_11054_40476# a_11054_40124# 0.010937f
C1322 XA0.XA1.XA1.MP3.G a_n178_39420# 0.023111f
C1323 XA3.XA1.CHL_OP D<5> 0.208613f
C1324 XA8.XA1.CHL_OP AVDD 2.05768f
C1325 XA6.XA6.Y XA6.XA8.A 0.527529f
C1326 a_11054_2446# a_11054_2094# 0.010937f
C1327 XB1.XA1.Y XB1.XA1.MP0.G 0.22339f
C1328 XA0.CEO XA0.XA11.Y 0.158152f
C1329 a_11054_44348# XA4.CN1 0.066018f
C1330 XA4.XA1.CHL_OP a_9902_43468# 0.010411f
C1331 a_9614_686# CK_SAMPLE_BSSW 0.071059f
C1332 XDAC2.XC128a<1>.XRES16.B D<8> 0.031495f
C1333 XB1.TIE_L SAR_IN 0.542565f
C1334 XA8.XA10.Y AVDD 0.721072f
C1335 XA2.XA10.Y VREF 0.011196f
C1336 XA2.XA1.XA4.LCK_N XA2.XA1.XA4.MN1.S 0.030434f
C1337 XA3.XA10.A XA3.XA8.A 0.062692f
C1338 XA0.XA1.XA1.MP3.S a_974_40476# 0.04865f
C1339 a_13574_40828# a_13574_40476# 0.010937f
C1340 XA5.XA6.MN1.S CK_SAMPLE 0.053284f
C1341 XA4.CN0 D<1> 0.073242f
C1342 a_18614_39420# a_18614_39068# 0.010937f
C1343 a_17462_41884# AVDD 0.397775f
C1344 a_19982_47340# a_19982_46988# 0.010937f
C1345 XA4.ENO a_11054_46988# 0.077282f
C1346 a_n178_41884# EN 0.076552f
C1347 XDAC2.XC0.XRES16.B XDAC2.XC0.XRES1A.B 0.467299f
C1348 a_8462_2974# AVDD 0.471212f
C1349 XB1.XA4.GNG m3_7598_2200# 0.105547f
C1350 XA6.CP0 XA6.XA1.CHL_OP 0.729561f
C1351 a_974_45228# XA0.XA1.CHL_OP 0.066018f
C1352 XA4.EN XA3.XA1.XA4.LCK_N 0.154232f
C1353 XA0.ENO a_2342_39420# 0.01235f
C1354 SAR_IP CK_SAMPLE_BSSW 0.016648f
C1355 a_16094_47340# AVDD 0.390024f
C1356 XA0.CMP_OP D<1> 0.072437f
C1357 XA8.XA2.A VREF 0.384473f
C1358 XA6.XA2.A EN 0.166272f
C1359 XA5.ENO XA5.CN1 0.083825f
C1360 XA8.XA11.Y XA8.XA11.MP1.S 0.054448f
C1361 a_19982_43468# XA8.XA2.A 0.067588f
C1362 XA7.ENO XA7.XA1.XA1.MP3.S 0.077008f
C1363 XDAC1.X16ab.XRES8.B SARP 27.705599f
C1364 XDAC2.XC1.XRES16.B SARN 55.2953f
C1365 XA0.CMP_OP XA0.XA1.XA1.MN2.S 0.024478f
C1366 XA0.CMP_ON a_14942_40124# 0.074163f
C1367 XA4.XA1.XA1.MP3.G a_11054_39772# 0.033843f
C1368 XA7.XA1.CHL_OP AVDD 2.02278f
C1369 a_21134_45228# D<0> 0.017384f
C1370 XA6.XA6.Y XA6.XA9.MN1.S 0.023798f
C1371 a_9614_2270# XB1.XA1.MP0.G 0.098163f
C1372 XA0.CN0 XA5.CN0 0.172071f
C1373 XA1.CN0 XA4.CN0 0.153041f
C1374 XA2.CN0 XA3.CN0 2.0007f
C1375 a_n178_49452# a_n178_49100# 0.010937f
C1376 a_11054_49452# XA4.XA11.Y 0.066018f
C1377 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES8.B 0.477132f
C1378 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES2.B 0.015267f
C1379 a_8462_686# CK_SAMPLE_BSSW 0.067588f
C1380 a_9902_44348# XA4.CN1 0.069545f
C1381 XA4.ENO XA5.XA1.XA4.MN2.S 0.012065f
C1382 a_11054_686# SAR_IP 0.060109f
C1383 XDAC2.XC1.XRES8.B XDAC2.XC1.XRES2.B 0.446669f
C1384 XB1.TIE_L SAR_IP 0.537987f
C1385 XA7.XA10.Y AVDD 0.714772f
C1386 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES16.B 0.063821f
C1387 XA1.XA10.Y VREF 0.01109f
C1388 XA0.CMP_OP a_4862_41180# 0.085247f
C1389 XA3.XA10.A XA3.XA6.Y 0.205884f
C1390 XA0.XA1.XA1.MP3.G a_974_40476# 0.098305f
C1391 XA3.CN0 SARP 0.032152f
C1392 XA4.CN0 D<2> 0.066013f
C1393 XA4.XA6.MP1.S D<4> 0.016737f
C1394 XA5.XA6.MP1.S CK_SAMPLE 0.022628f
C1395 a_16094_41884# AVDD 0.397775f
C1396 XA4.ENO a_9902_46988# 0.066245f
C1397 XA1.XA6.Y XA1.CP0 0.010942f
C1398 XA8.XA6.Y XA8.XA6.MP1.S 0.055045f
C1399 XA1.CN0 XA0.CMP_OP 0.055878f
C1400 XB1.XA4.GNG m3_7526_2200# 0.0666f
C1401 XA7.CN0 XA0.CMP_ON 0.061266f
C1402 a_n178_45228# XA0.XA1.CHL_OP 0.06825f
C1403 XA2.ENO XA3.XA1.XA4.LCK_N 0.3401f
C1404 XA4.EN XA4.XA1.XA5.MN2.S 0.010423f
C1405 a_21134_49804# AVDD 0.450198f
C1406 XDAC2.XC32a<0>.XRES1A.B XDAC2.XC64a<0>.XRES1B.B 0.62895f
C1407 a_6014_48572# XA2.XA10.A 0.066018f
C1408 XA0.ENO a_974_39420# 0.010025f
C1409 XA6.ENO a_16094_39772# 0.054233f
C1410 XA8.XA1.CHL_OP XA8.XA1.XA4.MN2.S 0.062799f
C1411 XA1.XA1.XA5.MN2.S XA1.XA1.XA5.MN1.S 0.050207f
C1412 SAR_IP SAR_IN 0.010593f
C1413 a_3494_41180# a_3494_40828# 0.010937f
C1414 a_19982_40124# a_19982_39772# 0.010937f
C1415 XA7.XA2.A VREF 0.387511f
C1416 XA0.CMP_OP D<2> 0.071274f
C1417 a_12422_47692# a_12422_47340# 0.010937f
C1418 XA5.XA2.A EN 0.166192f
C1419 a_12422_1038# a_12422_686# 0.010937f
C1420 XA7.XA1.XA1.MN2.S D<1> 0.023009f
C1421 a_7382_40124# AVDD 0.3588f
C1422 XDAC1.XC128a<1>.XRES8.B XDAC1.XC128a<1>.XRES16.B 0.1057f
C1423 XA8.XA11.Y XA8.XA10.Y 0.098057f
C1424 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES1A.B 0.022835f
C1425 XA6.XA1.CHL_OP XA6.XA1.XA5.MN2.S 0.013533f
C1426 XA5.XA1.CHL_OP XA5.XA1.XA4.LCK_N 0.204048f
C1427 XA7.ENO XA7.XA1.XA1.MP3.G 0.316693f
C1428 XA1.ENO a_2342_40476# 0.016912f
C1429 XDAC1.XC1.XRES2.B SARP 7.01088f
C1430 XA0.CMP_ON a_13574_40124# 0.072592f
C1431 XA3.XA1.XA4.MP2.S XA3.XA1.XA4.MP1.S 0.050207f
C1432 a_9902_40476# a_9902_40124# 0.010937f
C1433 XA6.XA1.CHL_OP AVDD 2.02306f
C1434 a_17462_45228# VREF 0.059568f
C1435 XA2.XA1.CHL_OP D<6> 0.208852f
C1436 XA1.XA8.A a_3494_47692# 0.160931f
C1437 a_8462_2270# XB1.XA1.MP0.G 0.067588f
C1438 a_9614_2270# XB1.XA1.Y 0.015779f
C1439 a_12422_40828# AVDD 0.407021f
C1440 XA2.CN0 XA2.XA6.MP1.S 0.028026f
C1441 a_17462_41180# EN 0.072753f
C1442 a_9902_49452# XA4.XA11.Y 0.070936f
C1443 a_11054_49452# XA4.CEO 0.040807f
C1444 XA3.XA1.CHL_OP a_8534_43468# 0.010411f
C1445 a_15014_n18# AVDD 0.44936f
C1446 a_11054_686# SARP 0.038089f
C1447 XDAC2.XC128a<1>.XRES16.B SARN 55.2956f
C1448 XB1.TIE_L SARP 0.561505f
C1449 XA7.XA11.MP1.S AVDD 0.101676f
C1450 XA8.XA1.XA5.MP2.S XA8.XA1.XA5.MP1.S 0.050207f
C1451 XA5.XA1.XA4.LCK_N a_13574_41884# 0.031412f
C1452 XA2.CN1 XA2.XA1.XA1.MP3.G 0.012171f
C1453 XA0.CMP_OP a_3494_41180# 0.086948f
C1454 XA0.XA1.XA1.MP3.G a_n178_40476# 0.066018f
C1455 a_12422_40828# a_12422_40476# 0.010937f
C1456 XA4.CN0 D<3> 0.097821f
C1457 XA3.CN0 EN 0.064814f
C1458 a_17462_39420# a_17462_39068# 0.010937f
C1459 XA4.XA6.Y a_11054_46108# 0.023316f
C1460 a_18614_47340# a_18614_46988# 0.010937f
C1461 XA8.XA6.Y XA8.XA6.MN1.S 0.026506f
C1462 XDAC1.XC0.XRES16.B XDAC1.XC0.XRES1A.B 0.467299f
C1463 a_8462_3326# AVDD 0.45186f
C1464 XB1.XA4.GNG m3_974_3000# 0.024512f
C1465 XA5.CP0 XA5.XA1.CHL_OP 0.729665f
C1466 a_4862_48572# XA2.XA10.A 0.068275f
C1467 XA8.XA2.A XA8.XA1.XA5.MN2.S 0.050207f
C1468 SARP SAR_IN 0.696352f
C1469 XA6.XA2.A VREF 0.387511f
C1470 XA0.CMP_OP D<3> 0.072437f
C1471 XA7.XA8.A XA7.ENO 0.144331f
C1472 XA4.XA2.A EN 0.166272f
C1473 a_7382_42588# AVDD 0.376544f
C1474 XB1.XA3.B a_8462_334# 0.011407f
C1475 XB2.XA3.MP0.S a_15014_686# 0.023111f
C1476 XA4.ENO XA4.CN1 0.083825f
C1477 XA0.CN0 XA0.XA1.CHL_OP 0.036653f
C1478 a_6014_40124# AVDD 0.358987f
C1479 a_18614_43468# XA7.XA2.A 0.066018f
C1480 XA6.ENO XA7.XA1.XA1.MP3.G 0.126806f
C1481 XA0.CMP_OP a_21134_40476# 0.067407f
C1482 XA0.CMP_ON a_12422_40124# 0.067588f
C1483 XA8.XA1.XA1.MP3.G a_21134_40124# 0.028807f
C1484 XA5.XA1.CHL_OP AVDD 2.02278f
C1485 a_16094_45228# VREF 0.059568f
C1486 XA1.XA6.Y a_3494_47692# 0.017683f
C1487 XA1.XA8.A a_2342_47692# 0.133834f
C1488 a_8462_2270# XB1.XA1.Y 0.030771f
C1489 a_15014_2622# a_15014_2270# 0.010937f
C1490 a_11054_40828# AVDD 0.407021f
C1491 a_16094_41180# EN 0.074323f
C1492 a_9902_49452# XA4.CEO 0.023111f
C1493 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES8.B 0.029725f
C1494 XDAC2.XC64b<1>.XRES16.B XDAC2.X16ab.XRES16.B 0.010386f
C1495 a_8534_44348# XA3.CN1 0.067974f
C1496 a_12422_1038# SAR_IN 0.067687f
C1497 XA20.XA2.N1 XA0.CMP_ON 0.114494f
C1498 XDAC1.XC128a<1>.XRES2.B SARP 7.01089f
C1499 XDAC1.XC1.XRES8.B XDAC1.XC1.XRES2.B 0.446669f
C1500 XA6.XA11.MP1.S AVDD 0.118921f
C1501 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES16.B 0.063821f
C1502 XA2.XA10.A XA2.XA8.A 0.062692f
C1503 XA4.XA1.XA1.MP3.G XA4.XA1.XA1.MP3.S 0.073693f
C1504 XA2.CN1 XDAC2.XC32a<0>.XRES16.B 0.018765f
C1505 XA5.XA6.MP1.S AVDD 0.092671f
C1506 XA3.CN0 D<8> 0.173434f
C1507 XA4.CN0 D<4> 1.79262f
C1508 XA4.EN a_8534_46988# 0.067815f
C1509 XA8.XA1.XA5.MP1.S EN 0.030477f
C1510 XA8.XA6.Y XA8.CN0 0.093605f
C1511 XB1.XA4.GNG m3_830_3000# 0.049023f
C1512 XA2.ENO XA3.XA1.XA5.MN2.S 0.010423f
C1513 XA2.CN0 XA2.XA2.A 0.028f
C1514 a_23654_45404# XA20.XA2.VMR 0.023111f
C1515 XA20.XA1.CKN a_23654_39420# 0.070731f
C1516 XA5.ENO a_14942_39772# 0.085451f
C1517 XA7.XA1.CHL_OP XA7.XA1.XA4.MN2.S 0.062799f
C1518 XA0.CMP_ON a_19982_41884# 0.087868f
C1519 XA1.XA1.XA5.MN2.S XA1.XA1.XA4.LCK_N 0.010898f
C1520 SARP SAR_IP 0.997754f
C1521 a_2342_41180# a_2342_40828# 0.010937f
C1522 XA20.XA1.CKN SARN 0.904997f
C1523 a_12422_47340# AVDD 0.390024f
C1524 a_18614_40124# a_18614_39772# 0.010937f
C1525 a_23654_47692# XA20.XA1.CKN 0.031543f
C1526 XA5.XA2.A VREF 0.387511f
C1527 a_11054_47692# a_11054_47340# 0.010937f
C1528 XA3.XA6.Y a_8534_46988# 0.047651f
C1529 XA7.XA6.Y XA7.ENO 0.051732f
C1530 XA0.CMP_OP D<4> 0.071274f
C1531 XA3.XA2.A EN 0.166192f
C1532 a_6014_42588# AVDD 0.376544f
C1533 a_11054_1038# a_11054_686# 0.010937f
C1534 XB2.XA3.MP0.S a_13862_686# 0.036577f
C1535 XA7.CEO XA8.XA11.MP1.S 0.010771f
C1536 XDAC2.XC128a<1>.XRES8.B XDAC2.XC128a<1>.XRES2.B 0.446669f
C1537 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES16.B 0.063821f
C1538 XA5.XA1.CHL_OP XA5.XA1.XA5.MN2.S 0.013533f
C1539 XDAC2.X16ab.XRES8.B SARN 27.705599f
C1540 a_17462_43468# XA7.XA2.A 0.067827f
C1541 XA0.ENO a_974_40476# 0.017441f
C1542 XA6.ENO XA6.XA1.XA1.MP3.S 0.076247f
C1543 XA0.CMP_OP a_19982_40476# 0.090364f
C1544 XA0.CMP_ON a_11054_40124# 0.066018f
C1545 XA7.XA1.XA4.LCK_N a_18614_41180# 0.060353f
C1546 a_8534_40476# a_8534_40124# 0.010937f
C1547 XA4.XA1.CHL_OP AVDD 2.02306f
C1548 XA1.XA1.CHL_OP D<7> 0.208613f
C1549 XA0.CN0 XA4.CN0 0.172401f
C1550 a_7382_44348# XA3.CN1 0.067588f
C1551 XA20.XA2.N1 a_23654_43996# 0.035229f
C1552 XB2.XA3.B CK_SAMPLE_BSSW 0.059546f
C1553 XA6.XA10.Y AVDD 0.717498f
C1554 XA0.XA10.Y VREF 0.011196f
C1555 XA8.XA1.XA4.LCK_N XA8.XA1.XA5.MN1.S 0.030434f
C1556 XA2.XA10.A XA2.XA9.MN1.S 0.073313f
C1557 a_11054_40828# a_11054_40476# 0.010937f
C1558 XA7.XA6.MP3.S AVDD 0.112857f
C1559 XA2.CN0 SARP 0.03275f
C1560 XA3.CN0 VREF 0.49936f
C1561 XA5.CN0 CK_SAMPLE 0.075434f
C1562 a_16094_39420# a_16094_39068# 0.010937f
C1563 a_12422_41884# AVDD 0.397775f
C1564 a_17462_47340# a_17462_46988# 0.010937f
C1565 XA4.EN a_7382_46988# 0.075712f
C1566 a_23654_47164# XA20.XA1.CK 0.036577f
C1567 XDAC2.XC0.XRES2.B XDAC2.XC0.XRES1A.B 0.015267f
C1568 XA0.CN0 XA0.CMP_OP 0.057021f
C1569 XB1.XA4.GNG m3_7598_3160# 0.105547f
C1570 a_22502_39068# AVDD 0.442014f
C1571 XA6.CN0 XA0.CMP_ON 0.062575f
C1572 a_23654_45404# XA20.XA2.CO 0.066018f
C1573 XA4.CP0 XA4.XA1.CHL_OP 0.729561f
C1574 a_3494_48572# XA1.XA10.A 0.066704f
C1575 XA8.XA10.Y XA8.XA10.A 0.201839f
C1576 a_17462_49804# AVDD 0.451537f
C1577 XDAC1.XC32a<0>.XRES1A.B XDAC1.XC64a<0>.XRES1B.B 0.62895f
C1578 XA20.XA1.CKN a_22502_39420# 0.066018f
C1579 XA7.XA2.A XA7.XA1.XA5.MN2.S 0.050207f
C1580 XA0.CMP_ON a_18614_41884# 0.095246f
C1581 XA4.CEIN XA3.XA6.Y 0.021942f
C1582 VREF CK_SAMPLE_BSSW 0.045361f
C1583 a_11054_47340# AVDD 0.390024f
C1584 XA7.XA2.A D<1> 0.040084f
C1585 XA4.XA2.A VREF 0.387511f
C1586 XA3.XA6.Y a_7382_46988# 0.023982f
C1587 XA2.XA2.A EN 0.166272f
C1588 XA0.CMP_OP D<5> 0.063761f
C1589 XA4.EN XA3.CN1 0.195951f
C1590 XA7.CN0 a_17462_46108# 0.101833f
C1591 XA7.CEO XA8.XA10.Y 0.303978f
C1592 XA7.XA11.Y XA7.XA10.Y 0.098057f
C1593 XDAC1.X16ab.XRES4.B SARP 13.9307f
C1594 XA6.ENO XA6.XA1.XA1.MP3.G 0.363295f
C1595 XDAC2.XC1.XRES2.B SARN 7.01088f
C1596 XA0.XA6.Y VREF 0.078171f
C1597 XA0.CMP_OP a_18614_40476# 0.088673f
C1598 XA0.CMP_ON a_9902_40124# 0.074163f
C1599 XA7.XA1.XA4.LCK_N a_17462_41180# 0.023475f
C1600 XA0.XA6.Y XA0.DONE 0.014904f
C1601 XA5.XA8.A XA5.XA9.MN1.S 0.010335f
C1602 XA5.XA6.Y XA6.XA6.Y 0.046858f
C1603 XA3.XA1.CHL_OP AVDD 2.02278f
C1604 a_17462_45228# D<1> 0.017384f
C1605 a_13862_2622# a_13862_2270# 0.010937f
C1606 a_8534_49452# XA3.XA11.Y 0.069366f
C1607 XDAC1.XC64b<1>.XRES16.B XDAC1.X16ab.XRES16.B 0.010386f
C1608 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES8.B 0.029725f
C1609 XA20.XA2.N1 a_22502_43996# 0.023357f
C1610 XB2.XA3.B SAR_IN 0.241597f
C1611 a_11054_1038# SAR_IP 0.067687f
C1612 a_12422_686# SARN 0.037937f
C1613 XA8.XA1.CHL_OP XA0.CMP_ON 0.161448f
C1614 XA5.CN0 XA5.XA1.XA4.LCK_N 0.01537f
C1615 XA5.XA10.Y AVDD 0.714772f
C1616 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES16.B 0.05157f
C1617 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES2.B 0.033713f
C1618 XB1.TIE_L VREF 0.057694f
C1619 XA2.XA1.XA4.LCK_N XA2.XA1.XA4.MN2.S 0.030434f
C1620 XA1.CN1 XA1.XA1.XA1.MP3.G 0.012023f
C1621 XA0.CMP_OP a_n178_41180# 0.085247f
C1622 XA2.XA10.A XA2.XA6.Y 0.205884f
C1623 XA6.XA6.MP3.S AVDD 0.112857f
C1624 XA3.CN0 SARN 0.048999f
C1625 XA4.XA6.MP1.S CK_SAMPLE 0.022425f
C1626 XA2.CN0 EN 0.065579f
C1627 a_11054_41884# AVDD 0.397775f
C1628 XA8.XA1.XA5.MP2.S EN 0.044228f
C1629 a_22502_47164# XA20.XA1.CK 0.023111f
C1630 XB1.XA4.GNG m3_7526_3160# 0.0666f
C1631 XA7.CN0 XA7.CN1 0.050499f
C1632 a_21134_39068# AVDD 0.443169f
C1633 XB2.XA4.GNG XDAC2.XC1.XRES1A.B 0.403704f
C1634 a_22502_45404# XA20.XA2.CO 0.067974f
C1635 a_2342_48572# XA1.XA10.A 0.067588f
C1636 a_16094_49804# AVDD 0.450382f
C1637 XA0.CMP_ON a_17462_41884# 0.011704f
C1638 XA1.XA1.XA5.MP2.S XA1.XA1.XA5.MP1.S 0.050207f
C1639 XA4.ENO a_13574_39772# 0.082231f
C1640 XA5.ENO a_12422_39772# 0.044989f
C1641 XA0.CMP_OP XA6.XA1.XA4.LCK_N 0.375196f
C1642 a_974_41180# a_974_40828# 0.010937f
C1643 a_17462_40124# a_17462_39772# 0.010937f
C1644 a_9902_47692# a_9902_47340# 0.010937f
C1645 XA6.XA8.A XA6.ENO 0.144331f
C1646 XA0.CMP_OP D<6> 0.062543f
C1647 XA3.XA2.A VREF 0.387511f
C1648 XA1.XA2.A EN 0.166192f
C1649 XA6.XA1.XA1.MN2.S D<2> 0.026904f
C1650 XA2.ENO XA3.CN1 0.239401f
C1651 XA5.CN0 XA5.CP0 0.796454f
C1652 a_2342_40124# AVDD 0.3588f
C1653 XA7.XA11.Y XA7.XA11.MP1.S 0.054448f
C1654 XA7.CEO XA7.XA10.Y 0.13078f
C1655 XDAC1.XC128a<1>.XRES8.B XDAC1.XC128a<1>.XRES2.B 0.446669f
C1656 XDAC2.XC128b<2>.XRES2.B XDAC2.XC128b<2>.XRES16.B 0.470901f
C1657 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES16.B 0.063821f
C1658 a_16094_43468# XA6.XA2.A 0.066256f
C1659 XA5.ENO XA6.XA1.XA1.MP3.G 0.031841f
C1660 XDAC1.XC1.XRES8.B SARP 27.705599f
C1661 XA2.XA1.XA4.MP2.S XA2.XA1.XA4.MP1.S 0.050207f
C1662 XA0.CMP_OP a_17462_40476# 0.068716f
C1663 XA0.CMP_ON a_8534_40124# 0.072592f
C1664 XA3.XA1.XA1.MP3.G a_7382_39772# 0.033843f
C1665 a_7382_40476# a_7382_40124# 0.010937f
C1666 XA5.XA6.Y XA5.XA9.MN1.S 0.023798f
C1667 XA0.XA8.A a_974_47692# 0.133834f
C1668 XA2.XA1.CHL_OP AVDD 2.02306f
C1669 a_12422_45228# VREF 0.059568f
C1670 XB2.XA2.MP0.G XB2.XA1.MP0.G 0.010347f
C1671 a_7382_40828# AVDD 0.407021f
C1672 a_12422_41180# EN 0.072753f
C1673 a_8534_49452# XA4.CEIN 0.024074f
C1674 a_7382_49452# XA3.XA11.Y 0.067588f
C1675 a_6014_44348# XA2.CN1 0.066018f
C1676 XA2.XA1.CHL_OP a_4862_43468# 0.010411f
C1677 XB1.XA3.B CK_SAMPLE_BSSW 0.059546f
C1678 a_11054_1038# SARP 0.045536f
C1679 XB2.XA3.MP0.S SAR_IN 0.100365f
C1680 XA7.XA1.CHL_OP XA0.CMP_ON 0.305949f
C1681 XDAC2.XC128a<1>.XRES2.B SARN 7.01089f
C1682 XB1.TIE_L SARN 0.390145f
C1683 XA5.XA11.MP1.S AVDD 0.101676f
C1684 XA1.XA1.XA4.LCK_N XA1.XA1.XA4.MN1.S 0.030434f
C1685 XA0.CMP_OP XA8.XA1.XA4.MP1.S 0.026047f
C1686 a_9902_40828# a_9902_40476# 0.010937f
C1687 XA5.CN0 AVDD 4.50659f
C1688 XA2.CN0 D<8> 0.179097f
C1689 XA4.XA6.MN1.S CK_SAMPLE 0.050648f
C1690 a_14942_39420# a_14942_39068# 0.010937f
C1691 a_16094_47340# a_16094_46988# 0.010937f
C1692 XA8.ENO XA20.XA1.CK 0.02089f
C1693 XA2.ENO a_6014_46988# 0.077282f
C1694 XA8.XA1.XA4.LCK_N EN 0.038188f
C1695 XDAC1.XC0.XRES2.B XDAC1.XC0.XRES1A.B 0.015267f
C1696 XB1.XA4.GNG m3_974_3960# 0.024512f
C1697 XA3.CP0 XA3.XA1.CHL_OP 0.745279f
C1698 XA7.XA10.Y XA7.XA10.A 0.201839f
C1699 XA0.CMP_ON a_16094_41884# 0.011248f
C1700 XA7.XA1.CHL_OP XA7.XA1.XA4.MP2.S 0.050207f
C1701 D<8> SARP 0.204103f
C1702 SARN SAR_IN 0.991833f
C1703 XA0.CN0 XDAC2.XC1.XRES16.B 0.028741f
C1704 XA8.XA8.A a_21134_47340# 0.091063f
C1705 XA0.CMP_OP D<7> 0.063761f
C1706 XA2.XA2.A VREF 0.387511f
C1707 XA6.XA2.A D<2> 0.039281f
C1708 a_2342_42588# AVDD 0.376544f
C1709 XA0.XA2.A EN 0.206912f
C1710 XA2.ENO XA2.CN1 0.10108f
C1711 a_974_40124# AVDD 0.358987f
C1712 XA7.CEO XA7.XA11.MP1.S 0.012048f
C1713 XA4.XA1.CHL_OP XA4.XA1.XA5.MN1.S 0.011494f
C1714 XA20.XA1.CKN XA20.XA1.MP0.S 0.109021f
C1715 XA5.ENO XA5.XA1.XA1.MP3.S 0.077008f
C1716 a_14942_43468# XA6.XA2.A 0.067588f
C1717 XA0.CMP_OP a_16094_40476# 0.067146f
C1718 XA0.CMP_ON a_7382_40124# 0.067588f
C1719 XA0.XA8.A a_n178_47692# 0.160931f
C1720 XA5.XA6.Y XA5.XA8.A 0.527529f
C1721 XA1.XA1.CHL_OP AVDD 2.02278f
C1722 a_11054_45228# VREF 0.059568f
C1723 a_16094_45228# D<2> 0.017384f
C1724 a_974_49804# AVDD 0.450382f
C1725 XA20.XA1.CK XA20.XA4.MP0.S 0.021464f
C1726 a_6014_40828# AVDD 0.407021f
C1727 a_11054_41180# EN 0.074323f
C1728 a_7382_49452# XA4.CEIN 0.029627f
C1729 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES4.B 0.430615f
C1730 a_4862_44348# XA2.CN1 0.069545f
C1731 a_8462_n18# AVDD 0.448205f
C1732 XA6.XA1.CHL_OP XA0.CMP_ON 0.231927f
C1733 XDAC1.XC128a<1>.XRES8.B SARP 27.705599f
C1734 XA4.XA11.MP1.S AVDD 0.118921f
C1735 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES16.B 0.05157f
C1736 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES2.B 0.033713f
C1737 XA0.CMP_OP XA8.XA1.XA4.MN1.S 0.036081f
C1738 XA1.XA10.A XA1.XA9.MN1.S 0.073313f
C1739 XA3.XA1.XA1.MP3.G XA3.XA1.XA1.MP3.S 0.073693f
C1740 a_21134_40828# XA8.XA1.XA1.MP3.G 0.069927f
C1741 XA4.XA6.MP1.S AVDD 0.092671f
C1742 XA3.CN0 D<1> 0.076653f
C1743 XA2.CN0 VREF 0.496795f
C1744 XA5.XA6.MP3.S D<3> 0.028396f
C1745 XA4.CN0 CK_SAMPLE 0.075021f
C1746 XA7.XA6.Y XA7.XA6.MN1.S 0.026506f
C1747 XA2.ENO a_4862_46988# 0.066245f
C1748 XB1.XA4.GNG m3_830_3960# 0.049023f
C1749 XA8.CP0 a_21134_45228# 0.070763f
C1750 a_974_48572# XA0.XA10.A 0.066018f
C1751 XA0.CMP_ON a_14942_41884# 0.090551f
C1752 XA4.ENO a_11054_39772# 0.054233f
C1753 XA7.XA2.A XA7.XA1.XA5.MP2.S 0.050207f
C1754 D<8> EN 0.339177f
C1755 SARN SAR_IP 0.806807f
C1756 a_n178_41180# a_n178_40828# 0.010937f
C1757 a_7382_47340# AVDD 0.390024f
C1758 a_16094_40124# a_16094_39772# 0.010937f
C1759 XA20.XA10.A XA20.XA10.MN1.S 0.036164f
C1760 XA8.XA8.A a_19982_47340# 0.127528f
C1761 a_8534_47692# a_8534_47340# 0.010937f
C1762 XA6.XA6.Y XA6.ENO 0.051732f
C1763 XA1.XA2.A VREF 0.387511f
C1764 XA0.XA2.A D<8> 0.748414f
C1765 a_974_42588# AVDD 0.376544f
C1766 XA1.ENO XA2.CN1 0.344545f
C1767 XA5.XA1.XA1.MN2.S D<3> 0.023009f
C1768 XA6.CEO XA7.XA10.Y 0.352238f
C1769 XDAC1.XC128b<2>.XRES2.B XDAC1.XC128b<2>.XRES16.B 0.470901f
C1770 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES2.B 0.033713f
C1771 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES16.B 0.05157f
C1772 XA5.ENO XA5.XA1.XA1.MP3.G 0.316693f
C1773 XDAC2.X16ab.XRES4.B SARN 13.9307f
C1774 XA0.CMP_OP a_14942_40476# 0.09022f
C1775 XA0.CMP_ON a_6014_40124# 0.066018f
C1776 XA7.XA1.XA1.MP3.G a_17462_40124# 0.028807f
C1777 a_6014_40476# a_6014_40124# 0.010937f
C1778 XA0.XA1.CHL_OP AVDD 2.02312f
C1779 XA1.CN0 XA3.CN0 0.15748f
C1780 XB1.XA3.B SAR_IP 0.241597f
C1781 XA1.XA1.CHL_OP a_3494_43468# 0.010411f
C1782 XA8.XA1.CHL_OP XA8.CN1 0.465167f
C1783 XA5.XA1.CHL_OP XA0.CMP_ON 0.30589f
C1784 a_15014_334# AVDD 0.490722f
C1785 XA4.XA10.Y AVDD 0.717498f
C1786 XA0.CMP_OP XA8.XA1.XA4.MP2.S 0.011502f
C1787 XA8.XA1.XA5.MN2.S XA8.XA1.XA5.MN1.S 0.050207f
C1788 XA1.XA10.A XA1.XA8.A 0.062692f
C1789 a_19982_40828# XA8.XA1.XA1.MP3.G 0.067588f
C1790 a_8534_40828# a_8534_40476# 0.010937f
C1791 XA2.CN0 SARN 0.063034f
C1792 XA3.CN0 D<2> 0.069299f
C1793 XA6.XA6.MN3.S CK_SAMPLE 0.028011f
C1794 XA3.XA6.MP1.S D<5> 0.016737f
C1795 a_13574_39420# a_13574_39068# 0.010937f
C1796 XA8.XA6.Y XA8.XA6.MP3.S 0.055045f
C1797 XA7.XA6.Y XA7.XA6.MP1.S 0.055045f
C1798 XA3.XA6.Y a_7382_46108# 0.023316f
C1799 a_14942_47340# a_14942_46988# 0.010937f
C1800 a_7382_41884# AVDD 0.397775f
C1801 XA7.XA1.XA5.MP1.S EN 0.03516f
C1802 XDAC2.XC0.XRES2.B XDAC2.XC0.XRES16.B 0.470901f
C1803 XDAC2.XC0.XRES8.B XDAC2.XC0.XRES1A.B 0.029729f
C1804 XA2.ENO XA2.XA1.XA4.LCK_N 0.152052f
C1805 XA8.CP0 a_19982_45228# 0.101124f
C1806 XA2.CP0 XA2.XA1.CHL_OP 0.74533f
C1807 XB1.XA4.GNG m3_7598_4120# 0.105547f
C1808 a_17462_39068# AVDD 0.442014f
C1809 a_n178_48572# XA0.XA10.A 0.068275f
C1810 a_12422_49804# AVDD 0.451537f
C1811 XA0.CMP_ON a_13574_41884# 0.095246f
C1812 XA6.XA1.CHL_OP XA6.XA1.XA4.MP2.S 0.050207f
C1813 XA0.CMP_OP XA5.XA1.XA4.LCK_N 0.383512f
C1814 VREF EN 1.0181f
C1815 SARN SARP 5.60111f
C1816 a_6014_47340# AVDD 0.390024f
C1817 a_18614_47692# XA7.DONE 0.023111f
C1818 XA2.XA6.Y a_6014_46988# 0.023982f
C1819 XA0.XA2.A VREF 0.387511f
C1820 XA5.XA2.A D<3> 0.040084f
C1821 XB1.XA3.MP0.S a_9614_686# 0.036577f
C1822 XA0.CP1 XA0.XA1.CHL_OP 0.208852f
C1823 XA6.CN0 a_16094_46108# 0.103403f
C1824 XA0.ENO XA2.CN1 0.025149f
C1825 XA1.ENO XA1.CN1 0.193039f
C1826 XA8.XA1.XA1.MP2.S AVDD 0.068158f
C1827 XA6.CEO XA7.XA11.MP1.S 0.033093f
C1828 XA6.XA11.Y XA6.XA11.MP1.S 0.054448f
C1829 XA4.ENO XA5.XA1.XA1.MP3.G 0.126806f
C1830 a_13574_43468# XA5.XA2.A 0.066018f
C1831 XDAC1.X16ab.XRES1B.B SARP 3.63755f
C1832 XDAC2.XC1.XRES8.B SARN 27.705599f
C1833 XA0.CMP_OP a_13574_40476# 0.088673f
C1834 XA0.CMP_ON a_4862_40124# 0.074163f
C1835 XA2.XA1.XA1.MP3.G a_6014_39772# 0.033843f
C1836 XA20.XA2.VMR AVDD 4.96345f
C1837 a_9614_2622# a_9614_2270# 0.010937f
C1838 XA20.XA1.CKN a_23654_45404# 0.074595f
C1839 a_6014_49452# XA2.XA11.Y 0.066018f
C1840 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES4.B 0.430615f
C1841 a_3494_44348# XA1.CN1 0.067974f
C1842 XA4.EN XA4.XA1.XA4.MN2.S 0.012065f
C1843 XA4.XA1.CHL_OP XA0.CMP_ON 0.231927f
C1844 a_12422_1038# SARN 0.049644f
C1845 XB1.XA3.MP0.S SAR_IP 0.100365f
C1846 a_15014_1390# SAR_IN 0.023111f
C1847 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES2.B 0.015267f
C1848 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES8.B 0.477132f
C1849 XA3.XA10.Y AVDD 0.714772f
C1850 XA1.XA1.XA4.LCK_N XA1.XA1.XA4.MN2.S 0.030434f
C1851 XA0.CMP_OP XA7.XA1.XA4.MN1.S 0.027953f
C1852 XA1.XA10.A XA1.XA6.Y 0.205884f
C1853 XA5.XA6.MN3.S CK_SAMPLE 0.028011f
C1854 XA4.CN0 AVDD 4.40297f
C1855 XA4.XA6.MP3.S D<4> 0.028396f
C1856 XA3.CN0 D<3> 0.128372f
C1857 XA1.ENO a_3494_46988# 0.067815f
C1858 a_6014_41884# AVDD 0.397775f
C1859 XA7.XA1.XA4.LCK_N EN 0.038188f
C1860 XA1.ENO XA2.XA1.XA4.LCK_N 0.339883f
C1861 XA7.CN0 XA3.CN1 0.07141f
C1862 XA6.CN0 XA6.CN1 0.050966f
C1863 XB1.XA4.GNG m3_7526_4120# 0.0666f
C1864 a_16094_39068# AVDD 0.443169f
C1865 XB2.XA4.GNG XDAC2.XC1.XRES16.B 0.098205f
C1866 a_11054_49804# AVDD 0.450382f
C1867 XDAC2.XC32a<0>.XRES16.B XDAC2.XC32a<0>.XRES1A.B 0.467299f
C1868 XA0.CMP_ON a_12422_41884# 0.011704f
C1869 XA4.EN a_9902_39772# 0.085451f
C1870 XA6.XA2.A XA6.XA1.XA5.MP2.S 0.050207f
C1871 VREF D<8> 0.618337f
C1872 XA0.XA6.Y XA0.XA6.MP1.S 0.055045f
C1873 a_14942_40124# a_14942_39772# 0.010937f
C1874 a_17462_47692# XA7.DONE 0.023111f
C1875 a_7382_47692# a_7382_47340# 0.010937f
C1876 XA2.XA6.Y a_4862_46988# 0.047651f
C1877 XA0.CMP_OP AVDD 8.58774f
C1878 a_21134_43468# VREF 0.062695f
C1879 XB2.M1.G a_12422_n18# 0.067406f
C1880 XB1.XA3.MP0.S a_8462_686# 0.023111f
C1881 XA4.CN0 XA4.CP0 0.800576f
C1882 XA0.ENO XA1.CN1 0.239401f
C1883 XA8.XA1.XA1.MN2.S AVDD 0.045375f
C1884 XA6.CEO XA6.XA11.MP1.S 0.010609f
C1885 XA6.XA11.Y XA6.XA10.Y 0.098057f
C1886 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128b<2>.XRES16.B 0.1057f
C1887 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES2.B 0.033713f
C1888 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES16.B 0.05157f
C1889 XA4.ENO XA4.XA1.XA1.MP3.S 0.076247f
C1890 XA4.XA1.CHL_OP XA4.XA1.XA4.LCK_N 0.204048f
C1891 a_12422_43468# XA5.XA2.A 0.067827f
C1892 XDAC1.XC1.XRES4.B SARP 13.9307f
C1893 XA2.XA1.XA4.MN2.S XA2.XA1.XA4.MN1.S 0.050207f
C1894 XA0.CMP_OP a_12422_40476# 0.068716f
C1895 XA0.CMP_ON a_3494_40124# 0.072592f
C1896 a_4862_40476# a_4862_40124# 0.010937f
C1897 XA20.XA2.CO AVDD 4.68634f
C1898 a_7382_45228# VREF 0.059568f
C1899 XA20.XA1.CKN a_22502_45404# 0.066018f
C1900 a_2342_40828# AVDD 0.407021f
C1901 a_7382_41180# EN 0.072753f
C1902 a_6014_49452# XA2.CEO 0.040807f
C1903 a_4862_49452# XA2.XA11.Y 0.070936f
C1904 a_2342_44348# XA1.CN1 0.067588f
C1905 XA7.XA1.CHL_OP XA7.CN1 0.465167f
C1906 XA3.XA1.CHL_OP XA0.CMP_ON 0.30589f
C1907 a_13862_1390# SAR_IN 0.043386f
C1908 XA3.XA11.MP1.S AVDD 0.101676f
C1909 XDAC2.XC128a<1>.XRES8.B SARN 27.705599f
C1910 XA0.CMP_OP XA7.XA1.XA4.MP1.S 0.0111f
C1911 XA8.XA1.XA5.MN2.S XA8.XA1.XA4.LCK_N 0.010898f
C1912 XA7.XA1.XA4.LCK_N XA7.XA1.XA5.MN1.S 0.030434f
C1913 a_7382_40828# a_7382_40476# 0.010937f
C1914 XA2.CP0 XDAC1.X16ab.XRES16.B 0.018342f
C1915 XA3.XA6.MN1.S CK_SAMPLE 0.053284f
C1916 XA2.CN0 D<1> 0.079819f
C1917 XA3.CN0 D<4> 0.077262f
C1918 a_12422_39420# a_12422_39068# 0.010937f
C1919 XA7.ENO XA8.ENO 0.01884f
C1920 a_13574_47340# a_13574_46988# 0.010937f
C1921 XA1.ENO a_2342_46988# 0.075712f
C1922 XA8.XA1.XA5.MN2.S EN 0.016689f
C1923 XDAC1.XC0.XRES2.B XDAC1.XC0.XRES16.B 0.470901f
C1924 XDAC1.XC0.XRES8.B XDAC1.XC0.XRES1A.B 0.029729f
C1925 XA0.CP1 XA0.CMP_OP 0.062543f
C1926 XA7.CN0 XA2.CN1 0.159556f
C1927 XA7.CP0 a_18614_45228# 0.102695f
C1928 XA1.CP0 XA1.XA1.CHL_OP 0.745279f
C1929 a_23654_48924# a_23654_48572# 0.010937f
C1930 XA6.XA10.Y XA6.XA10.A 0.201839f
C1931 XA7.CN0 XA7.XA1.XA1.MP3.G 0.016018f
C1932 XA0.CMP_ON a_11054_41884# 0.011248f
C1933 XA0.XA1.XA5.MP2.S XA0.XA1.XA5.MP1.S 0.050207f
C1934 SARN D<8> 0.350364f
C1935 D<1> SARP 0.050623f
C1936 XA0.XA6.Y XA0.XA6.MN1.S 0.026506f
C1937 XA5.XA8.A XA5.ENO 0.144331f
C1938 XA8.XA6.Y a_19982_47340# 0.011912f
C1939 XA4.XA2.A D<4> 0.039281f
C1940 XB2.XA3.MP0.S XB2.XA3.B 0.098737f
C1941 XB1.TIE_L a_12422_1390# 0.067979f
C1942 XA7.XA1.XA1.MN2.S AVDD 0.036807f
C1943 XA6.CEO XA6.XA10.Y 0.02121f
C1944 XA4.ENO XA4.XA1.XA1.MP3.G 0.363295f
C1945 XA0.CMP_OP a_11054_40476# 0.067146f
C1946 XA0.CMP_ON a_2342_40124# 0.067588f
C1947 XA6.XA1.XA1.MP3.G a_16094_40124# 0.028807f
C1948 XA4.XA9.MN1.S XA4.XA8.A 0.010335f
C1949 a_21134_45228# AVDD 0.377363f
C1950 a_6014_45228# VREF 0.059568f
C1951 a_12422_45228# D<3> 0.017384f
C1952 a_8462_2622# a_8462_2270# 0.010937f
C1953 XA0.CN0 XA3.CN0 0.163814f
C1954 XA1.CN0 XA2.CN0 2.67683f
C1955 a_974_40828# AVDD 0.407021f
C1956 a_6014_41180# EN 0.074323f
C1957 a_4862_49452# XA2.CEO 0.023111f
C1958 XA2.ENO XA3.XA1.XA4.MN2.S 0.012065f
C1959 XA2.XA1.CHL_OP XA0.CMP_ON 0.231927f
C1960 XA3.CP0 XA0.CMP_OP 0.060463f
C1961 a_12422_1390# SAR_IN 0.056243f
C1962 XA2.XA11.MP1.S AVDD 0.118921f
C1963 XDAC1.XC128a<1>.XRES4.B SARP 13.9307f
C1964 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES2.B 0.015267f
C1965 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES8.B 0.477132f
C1966 XA0.CMP_OP XA8.XA1.XA4.MN2.S 0.014099f
C1967 XA0.XA10.A XA0.XA8.A 0.062692f
C1968 XA2.XA1.XA1.MP3.G XA2.XA1.XA1.MP3.S 0.073693f
C1969 a_18614_40828# XA7.XA1.XA1.MP3.G 0.066018f
C1970 XA3.XA6.MP1.S CK_SAMPLE 0.022628f
C1971 XA2.CN0 D<2> 0.072968f
C1972 XA3.CN0 D<5> 0.537393f
C1973 XA1.CN0 SARP 0.033203f
C1974 XA7.XA1.XA5.MN2.S EN 0.016683f
C1975 XA5.CN0 XA0.CMP_ON 0.060347f
C1976 XA1.CN0 XA1.XA2.A 0.02751f
C1977 XA7.CN0 XA1.CN1 0.076884f
C1978 XA7.CP0 a_17462_45228# 0.069193f
C1979 a_21134_39420# EN 0.067588f
C1980 XA0.CMP_ON a_9902_41884# 0.090551f
C1981 XA2.ENO a_8534_39772# 0.082231f
C1982 XA4.EN a_7382_39772# 0.044989f
C1983 XA6.XA1.CHL_OP XA6.XA1.XA4.MN2.S 0.062799f
C1984 D<2> SARP 0.046527f
C1985 D<1> EN 0.072241f
C1986 a_2342_47340# AVDD 0.390024f
C1987 XA0.XA6.Y XA0.CN0 0.093605f
C1988 a_13574_40124# a_13574_39772# 0.010937f
C1989 XA5.XA6.Y XA5.ENO 0.051732f
C1990 a_16094_47692# XA6.DONE 0.023111f
C1991 a_6014_47692# a_6014_47340# 0.010937f
C1992 a_22502_43116# AVDD 0.42631f
C1993 XB1.TIE_L a_11054_1390# 0.06903f
C1994 XA7.XA1.XA1.MP2.S AVDD 0.066893f
C1995 XA4.XA1.XA1.MN2.S D<4> 0.026904f
C1996 XA0.XA1.XA1.MN2.S EN 0.023301f
C1997 XA20.XA1.MP0.S SARP 0.255572f
C1998 XA5.CEO XA6.XA11.MP1.S 0.010771f
C1999 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128b<2>.XRES16.B 0.1057f
C2000 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES2.B 0.015267f
C2001 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES8.B 0.477132f
C2002 XA4.EN XA4.XA1.XA1.MP3.G 0.031841f
C2003 XA3.XA1.CHL_OP XA3.XA1.XA5.MN1.S 0.011494f
C2004 a_11054_43468# XA4.XA2.A 0.066256f
C2005 XDAC2.X16ab.XRES1B.B SARN 3.63755f
C2006 XA0.CMP_OP a_9902_40476# 0.09022f
C2007 XA0.CMP_ON a_974_40124# 0.066018f
C2008 a_3494_40476# a_3494_40124# 0.010937f
C2009 XA4.XA6.Y XA4.XA8.A 0.527529f
C2010 XA2.CP0 XA0.CMP_OP 0.060601f
C2011 XA1.XA1.CHL_OP XA0.CMP_ON 0.30589f
C2012 XA0.XA1.CHL_OP a_n178_43468# 0.010411f
C2013 XA6.XA1.CHL_OP XA6.CN1 0.465167f
C2014 XA2.XA10.Y AVDD 0.717498f
C2015 XA4.XA1.XA4.LCK_N a_9902_41884# 0.031412f
C2016 XA0.CMP_OP XA7.XA1.XA4.MN2.S 0.026188f
C2017 XA7.XA1.XA5.MN2.S XA7.XA1.XA5.MN1.S 0.050207f
C2018 a_17462_40828# XA7.XA1.XA1.MP3.G 0.071498f
C2019 a_6014_40828# a_6014_40476# 0.010937f
C2020 XA1.CN0 EN 0.064814f
C2021 XA2.CN0 D<3> 0.26947f
C2022 a_11054_39420# a_11054_39068# 0.010937f
C2023 XA6.ENO XA7.ENO 1.2771f
C2024 XA2.XA6.Y a_6014_46108# 0.023316f
C2025 a_12422_47340# a_12422_46988# 0.010937f
C2026 XA7.XA6.Y XA7.CN0 0.093605f
C2027 XA0.ENO a_974_46988# 0.077282f
C2028 a_2342_41884# AVDD 0.397775f
C2029 XA6.XA1.XA5.MP1.S EN 0.03516f
C2030 XDAC2.XC0.XRES8.B XDAC2.XC0.XRES16.B 0.1057f
C2031 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES1A.B 0.022835f
C2032 XA1.ENO XA1.XA1.XA4.LCK_N 0.154232f
C2033 XA0.CP0 XA0.XA1.CHL_OP 0.74533f
C2034 XA6.CN0 XA3.CN1 0.067614f
C2035 a_12422_39068# AVDD 0.442014f
C2036 a_7382_49804# AVDD 0.451537f
C2037 a_22502_48924# a_22502_48572# 0.010937f
C2038 XA5.XA10.Y XA5.XA10.A 0.201839f
C2039 XDAC1.XC32a<0>.XRES16.B XDAC1.XC32a<0>.XRES1A.B 0.467299f
C2040 XA0.CMP_ON a_8534_41884# 0.095246f
C2041 XA0.XA1.XA4.LCK_N XA0.XA1.XA5.MN1.S 0.030434f
C2042 D<1> D<8> 0.077821f
C2043 D<3> SARP 0.049966f
C2044 D<0> VREF 1.50643f
C2045 D<2> EN 0.07152f
C2046 XA20.XA1.CKN CK_SAMPLE 0.052735f
C2047 a_974_47340# AVDD 0.390024f
C2048 a_14942_47692# XA6.DONE 0.023111f
C2049 XA8.XA2.A AVDD 2.08545f
C2050 a_17462_43468# VREF 0.062747f
C2051 XA3.XA2.A D<5> 0.03176f
C2052 XB2.CKN a_15014_686# 0.120042f
C2053 XA6.XA1.XA1.MP2.S AVDD 0.068123f
C2054 XA5.CEO XA6.XA10.Y 0.303978f
C2055 XA5.XA11.Y XA5.XA10.Y 0.098057f
C2056 XA4.EN XA3.XA1.XA1.MP3.S 0.077008f
C2057 XA20.XA1.CK a_23654_40828# 0.140127f
C2058 a_9902_43468# XA4.XA2.A 0.067588f
C2059 XDAC1.XC64b<1>.XRES1A.B SARP 3.63804f
C2060 XDAC2.XC1.XRES4.B SARN 13.9307f
C2061 XA6.XA1.XA4.LCK_N a_16094_41180# 0.023475f
C2062 XA0.CMP_OP a_8534_40476# 0.088673f
C2063 XA0.CMP_ON a_n178_40124# 0.074097f
C2064 a_11054_45228# D<4> 0.017384f
C2065 XA4.XA6.Y XA4.XA9.MN1.S 0.023798f
C2066 XA8.ENO XA8.CN0 0.036889f
C2067 XA20.XA1.CK a_23654_46812# 0.101495f
C2068 a_21134_41180# AVDD 0.395845f
C2069 a_3494_49452# XA1.XA11.Y 0.069366f
C2070 XA1.CP0 XA0.CMP_OP 0.060463f
C2071 XA0.XA1.CHL_OP XA0.CMP_ON 0.231927f
C2072 a_8462_334# AVDD 0.492296f
C2073 a_12422_1390# SARP 0.025743f
C2074 a_11054_1390# SAR_IP 0.056243f
C2075 XA1.XA10.Y AVDD 0.714772f
C2076 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES8.B 0.029725f
C2077 XDAC2.XC64a<0>.XRES16.B XDAC2.XC1.XRES16.B 0.010386f
C2078 XA0.CMP_OP XA6.XA1.XA4.MP1.S 0.010745f
C2079 XA1.CN0 D<8> 0.089176f
C2080 XA2.XA6.MP1.S D<6> 0.016737f
C2081 XA3.XA6.MP1.S AVDD 0.092671f
C2082 XA2.CN0 D<4> 0.070487f
C2083 XA8.XA6.Y XA8.XA6.MN3.S 0.089305f
C2084 XA0.ENO a_n178_46988# 0.066245f
C2085 a_974_41884# AVDD 0.397775f
C2086 XA1.ENO XA2.XA1.XA5.MN2.S 0.010423f
C2087 XA0.ENO XA1.XA1.XA4.LCK_N 0.3401f
C2088 XA6.CP0 a_16094_45228# 0.070763f
C2089 XA6.CN0 XA2.CN1 0.303277f
C2090 XB2.XA4.GNG XDAC2.XC1.XRES2.B 0.010278f
C2091 XB1.XA4.GNG XDAC1.XC1.XRES1A.B 0.403704f
C2092 a_11054_39068# AVDD 0.443169f
C2093 a_6014_49804# AVDD 0.450382f
C2094 XDAC2.XC32a<0>.XRES2.B XDAC2.XC32a<0>.XRES1A.B 0.015267f
C2095 XA0.CMP_ON a_7382_41884# 0.011704f
C2096 XA0.XA1.XA5.MN2.S XA0.XA1.XA5.MN1.S 0.050207f
C2097 XA2.ENO a_6014_39772# 0.054233f
C2098 XA8.ENO a_21134_40124# 0.024823f
C2099 XA5.XA1.CHL_OP XA5.XA1.XA4.MN2.S 0.062799f
C2100 D<1> VREF 1.51304f
C2101 D<2> D<8> 0.086175f
C2102 D<4> SARP 0.050608f
C2103 D<3> EN 0.072241f
C2104 a_12422_40124# a_12422_39772# 0.010937f
C2105 XA1.XA6.Y a_3494_46988# 0.047651f
C2106 XA4.XA8.A XA4.ENO 0.144331f
C2107 XA7.XA8.A a_18614_47340# 0.129098f
C2108 a_4862_47692# a_4862_47340# 0.010937f
C2109 XA7.XA2.A AVDD 2.0645f
C2110 a_16094_43468# VREF 0.062747f
C2111 XB2.CKN a_13862_686# 0.113134f
C2112 XB1.M1.G a_11054_n18# 0.068977f
C2113 a_12422_1390# a_12422_1038# 0.010937f
C2114 XA6.XA1.XA1.MN2.S AVDD 0.036807f
C2115 XA3.XA1.XA1.MN2.S D<5> 0.023009f
C2116 XA5.XA11.Y XA5.XA11.MP1.S 0.054448f
C2117 XA5.CEO XA5.XA10.Y 0.13078f
C2118 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128b<2>.XRES2.B 0.446669f
C2119 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES16.B 0.063821f
C2120 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES2.B 0.015267f
C2121 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES8.B 0.477132f
C2122 XA4.EN XA3.XA1.XA1.MP3.G 0.316693f
C2123 XA20.XA1.CK a_22502_40828# 0.066143f
C2124 XA4.XA1.CHL_OP XA4.XA1.XA5.MN2.S 0.013533f
C2125 XA3.XA1.CHL_OP XA3.XA1.XA4.LCK_N 0.204048f
C2126 XDAC1.XC1.XRES1B.B SARP 3.63755f
C2127 XA6.XA1.XA4.LCK_N a_14942_41180# 0.060353f
C2128 XA1.XA1.XA4.MN2.S XA1.XA1.XA4.MN1.S 0.050207f
C2129 XA0.CMP_OP a_7382_40476# 0.068716f
C2130 XA1.XA1.XA1.MP3.G a_2342_39772# 0.033843f
C2131 a_2342_40476# a_2342_40124# 0.010937f
C2132 a_17462_45228# AVDD 0.377363f
C2133 a_2342_45228# VREF 0.059568f
C2134 a_12422_2798# a_12422_2446# 0.010937f
C2135 XA0.CN0 XA2.CN0 0.168345f
C2136 a_23654_47164# a_23654_46812# 0.010937f
C2137 a_2342_41180# EN 0.072753f
C2138 a_3494_49452# XA1.CEO 0.024074f
C2139 a_2342_49452# XA1.XA11.Y 0.067588f
C2140 XA20.XA2.VMR XA0.CMP_ON 0.16762f
C2141 XA0.CP0 XA0.CMP_OP 0.060601f
C2142 XA5.XA1.CHL_OP XA5.CN1 0.465167f
C2143 a_15014_686# AVDD 0.380767f
C2144 a_11054_1390# SARP 0.016378f
C2145 a_9614_1390# SAR_IP 0.043386f
C2146 XA1.XA11.MP1.S AVDD 0.101676f
C2147 XDAC2.XC128a<1>.XRES4.B SARN 13.9307f
C2148 XA0.CMP_OP XA6.XA1.XA4.MN1.S 0.024389f
C2149 XA7.XA1.XA5.MN2.S XA7.XA1.XA4.LCK_N 0.010898f
C2150 a_4862_40828# a_4862_40476# 0.010937f
C2151 XA2.CN0 D<5> 0.055822f
C2152 XA1.CN0 VREF 0.49936f
C2153 XA3.CN0 CK_SAMPLE 0.075434f
C2154 XA5.XA6.MP3.S AVDD 0.112857f
C2155 XA0.CN0 SARP 0.033467f
C2156 a_9902_39420# a_9902_39068# 0.010937f
C2157 XA5.ENO XA6.ENO 0.026181f
C2158 a_11054_47340# a_11054_46988# 0.010937f
C2159 XA7.XA1.XA4.LCK_N D<1> 0.019067f
C2160 XA7.XA1.XA5.MP2.S EN 0.044153f
C2161 XDAC1.XC0.XRES8.B XDAC1.XC0.XRES16.B 0.1057f
C2162 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES1A.B 0.022835f
C2163 XA4.CN0 XA0.CMP_ON 0.062602f
C2164 XA6.CP0 a_14942_45228# 0.101124f
C2165 XA6.CN0 XA1.CN1 0.073042f
C2166 a_17462_39420# EN 0.066018f
C2167 XA0.CMP_ON a_6014_41884# 0.011248f
C2168 XA6.XA2.A XA6.XA1.XA5.MN2.S 0.050207f
C2169 XA1.CEO XA1.XA6.Y 0.021942f
C2170 D<2> VREF 1.51285f
C2171 D<3> D<8> 0.073443f
C2172 D<5> SARP 0.090991f
C2173 D<1> SARN 0.038745f
C2174 D<4> EN 0.07152f
C2175 XA20.XA1.CKN AVDD 2.13851f
C2176 XA1.XA6.Y a_2342_46988# 0.023982f
C2177 XA2.XA2.A D<6> 0.03087f
C2178 XA6.XA2.A AVDD 2.06492f
C2179 a_13574_47692# XA5.DONE 0.023111f
C2180 XA7.XA6.Y a_18614_47340# 0.011912f
C2181 XA7.XA8.A a_17462_47340# 0.089492f
C2182 XB1.XA3.MP0.S XB1.XA3.B 0.098737f
C2183 XA8.CN0 XA8.XA6.MP1.S 0.028026f
C2184 XA5.XA1.XA1.MN2.S AVDD 0.036807f
C2185 XA5.CEO XA5.XA11.MP1.S 0.012048f
C2186 XA2.ENO XA3.XA1.XA1.MP3.G 0.126806f
C2187 XA0.CMP_ON XA0.CMP_OP 8.514441f
C2188 a_8534_43468# XA3.XA2.A 0.066018f
C2189 XA0.XA6.Y CK_SAMPLE 0.178114f
C2190 XA0.CMP_OP a_6014_40476# 0.067146f
C2191 XA0.CMP_ON XA8.XA1.XA1.MN2.S 0.064851f
C2192 XA0.CP1 XDAC1.XC128a<1>.XRES16.B 0.031495f
C2193 a_16094_45228# AVDD 0.377363f
C2194 a_974_45228# VREF 0.059568f
C2195 XB2.XA2.MP0.G a_15014_2622# 0.073828f
C2196 XA1.CN0 XA1.XA6.MP1.S 0.028026f
C2197 a_974_41180# EN 0.074323f
C2198 a_2342_49452# XA1.CEO 0.029627f
C2199 XDAC2.XC64b<1>.XRES1A.B XDAC2.X16ab.XRES1B.B 0.62895f
C2200 XA20.XA2.CO XA0.CMP_ON 0.477413f
C2201 XA4.CN0 XA4.XA1.XA4.LCK_N 0.015589f
C2202 a_8462_1390# SAR_IP 0.023111f
C2203 XB2.CKN CK_SAMPLE_BSSW 0.169642f
C2204 XA0.XA11.MP1.S AVDD 0.118921f
C2205 XDAC1.XC128a<1>.XRES1B.B SARP 3.63755f
C2206 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES8.B 0.029725f
C2207 XDAC1.XC64a<0>.XRES16.B XDAC1.XC1.XRES16.B 0.010386f
C2208 XA0.CMP_OP XA7.XA1.XA4.MP2.S 0.026257f
C2209 a_16094_40828# XA6.XA1.XA1.MP3.G 0.069927f
C2210 XA1.XA1.XA1.MP3.G XA1.XA1.XA1.MP3.S 0.073693f
C2211 XA1.CN0 SARN 0.179546f
C2212 XA2.XA6.MP1.S CK_SAMPLE 0.022425f
C2213 XA0.CN0 EN 0.067256f
C2214 XA2.CN0 D<6> 0.476007f
C2215 XA4.XA6.MP3.S AVDD 0.112857f
C2216 XA6.XA1.XA5.MP2.S EN 0.044228f
C2217 XA0.CN0 XA0.XA2.A 0.028f
C2218 XA0.ENO XA1.XA1.XA5.MN2.S 0.010423f
C2219 a_16094_39420# EN 0.067588f
C2220 XA8.XA10.Y a_21134_48572# 0.091063f
C2221 XA0.CMP_ON a_4862_41884# 0.090551f
C2222 XA6.CN0 XA6.XA1.XA1.MP3.G 0.021358f
C2223 XA1.ENO a_4862_39772# 0.085451f
C2224 XA0.CMP_OP XA4.XA1.XA4.LCK_N 0.375196f
C2225 D<2> SARN 0.034649f
C2226 D<3> VREF 1.51304f
C2227 D<4> D<8> 0.073479f
C2228 D<5> EN 0.064847f
C2229 D<6> SARP 0.084597f
C2230 XA0.XA6.Y XA0.XA6.MP3.S 0.055045f
C2231 XA7.DONE AVDD 0.241164f
C2232 a_11054_40124# a_11054_39772# 0.010937f
C2233 XA4.XA6.Y XA4.ENO 0.051732f
C2234 XA5.XA2.A AVDD 2.0645f
C2235 a_12422_47692# XA5.DONE 0.023111f
C2236 a_3494_47692# a_3494_47340# 0.010937f
C2237 XB2.M1.G a_12422_334# 0.158066f
C2238 a_13862_1390# XB2.XA3.MP0.S 0.071276f
C2239 a_11054_1390# a_11054_1038# 0.010937f
C2240 XB1.TIE_L XB2.CKN 0.066812f
C2241 XA5.XA1.XA1.MP2.S AVDD 0.066893f
C2242 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES8.B 0.029725f
C2243 XA4.CEO XA5.XA10.Y 0.352238f
C2244 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128b<2>.XRES2.B 0.446669f
C2245 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES16.B 0.063821f
C2246 XA2.ENO XA2.XA1.XA1.MP3.S 0.076247f
C2247 XA3.XA1.CHL_OP XA3.XA1.XA5.MN2.S 0.013533f
C2248 a_7382_43468# XA3.XA2.A 0.067827f
C2249 XDAC2.XC64b<1>.XRES1A.B SARN 3.63804f
C2250 XA0.CMP_OP a_4862_40476# 0.09022f
C2251 XA0.CMP_ON XA7.XA1.XA1.MN2.S 0.064851f
C2252 XA5.XA1.XA1.MP3.G a_12422_40124# 0.028807f
C2253 a_974_40476# a_974_40124# 0.010937f
C2254 XB1.XA2.MP0.G XB1.XA1.MP0.G 0.010347f
C2255 a_11054_2798# a_11054_2446# 0.010937f
C2256 XB2.XA2.MP0.G a_13862_2622# 0.066018f
C2257 a_22502_47164# a_22502_46812# 0.010937f
C2258 a_17462_41180# AVDD 0.39588f
C2259 XA20.XA2.CO a_23654_43996# 0.066264f
C2260 XA20.XA1.CK XA20.XA2.N2 0.034212f
C2261 XA8.XA1.CHL_OP a_21134_44348# 0.06801f
C2262 XA20.XA2.VMR a_22502_43996# 0.010987f
C2263 XA4.XA1.CHL_OP XA4.CN1 0.465167f
C2264 XB2.CKN SAR_IN 0.175642f
C2265 XA0.XA10.Y AVDD 0.717512f
C2266 XA0.CMP_OP XA6.XA1.XA4.MP2.S 0.026117f
C2267 XA7.XA1.XA5.MP2.S XA7.XA1.XA5.MP1.S 0.050207f
C2268 XA3.XA1.XA4.LCK_N a_8534_41884# 0.031412f
C2269 a_3494_40828# a_3494_40476# 0.010937f
C2270 a_14942_40828# XA6.XA1.XA1.MP3.G 0.067588f
C2271 XA2.XA6.MN1.S CK_SAMPLE 0.050648f
C2272 XA3.CN0 AVDD 4.48784f
C2273 XA0.CN0 D<8> 5.74687f
C2274 a_8534_39420# a_8534_39068# 0.010937f
C2275 a_22502_42236# AVDD 0.430438f
C2276 XA4.ENO XA5.ENO 1.2771f
C2277 XA6.XA1.XA4.LCK_N EN 0.038188f
C2278 a_9902_47340# a_9902_46988# 0.010937f
C2279 XA6.XA6.Y XA6.XA6.MP1.S 0.055045f
C2280 XDAC2.XC0.XRES8.B XDAC2.XC0.XRES2.B 0.446669f
C2281 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES16.B 0.063821f
C2282 XA7.ENO a_19982_42588# 0.070731f
C2283 XA5.CP0 a_13574_45228# 0.102695f
C2284 a_7382_39068# AVDD 0.442014f
C2285 a_2342_49804# AVDD 0.451537f
C2286 XDAC1.XC32a<0>.XRES2.B XDAC1.XC32a<0>.XRES1A.B 0.015267f
C2287 XA8.XA10.Y a_19982_48572# 0.13253f
C2288 XA4.XA10.Y XA4.XA10.A 0.201839f
C2289 XA0.CMP_ON a_3494_41884# 0.095246f
C2290 XA7.ENO a_18614_40124# 0.010898f
C2291 XA0.XA1.XA5.MN2.S XA0.XA1.XA4.LCK_N 0.010898f
C2292 XA5.XA1.CHL_OP XA5.XA1.XA4.MP2.S 0.050207f
C2293 XA5.XA2.A XA5.XA1.XA5.MN2.S 0.050207f
C2294 AVDD CK_SAMPLE_BSSW 19.8405f
C2295 D<3> SARN 0.034649f
C2296 D<6> EN 0.064085f
C2297 D<4> VREF 1.51285f
C2298 D<5> D<8> 0.073541f
C2299 D<7> SARP 0.139285f
C2300 XA0.XA6.Y XA0.XA6.MN3.S 0.089305f
C2301 XA6.DONE AVDD 0.241164f
C2302 XA20.XA1.MP0.S a_22502_39420# 0.023111f
C2303 XA1.XA2.A D<7> 0.03176f
C2304 XA4.XA2.A AVDD 2.06492f
C2305 a_12422_43468# VREF 0.062747f
C2306 XA4.XA1.XA1.MP2.S AVDD 0.068123f
C2307 a_974_49100# XB1.TIE_L 0.066018f
C2308 XA4.XA11.Y XA4.XA11.MP1.S 0.054448f
C2309 XA4.CEO XA5.XA11.MP1.S 0.033093f
C2310 XA2.ENO XA2.XA1.XA1.MP3.G 0.363295f
C2311 XDAC1.XC64b<1>.XRES16.B SARP 55.2956f
C2312 a_23654_48220# DONE 0.066018f
C2313 XA0.XA6.Y AVDD 0.864427f
C2314 XDAC2.XC1.XRES1B.B SARN 3.63755f
C2315 XA0.CMP_OP a_3494_40476# 0.088673f
C2316 XA0.XA1.XA1.MP3.G a_974_39772# 0.033843f
C2317 XA3.XA8.A XA3.XA9.MN1.S 0.010335f
C2318 XA3.XA6.Y XA4.XA6.Y 0.046858f
C2319 a_7382_45228# D<5> 0.017384f
C2320 XA8.XA1.XA4.MP1.S EN 0.027192f
C2321 a_16094_41180# AVDD 0.39588f
C2322 a_974_49452# XA0.XA11.Y 0.066018f
C2323 XDAC1.XC64b<1>.XRES1A.B XDAC1.X16ab.XRES1B.B 0.62895f
C2324 XA8.XA1.CHL_OP a_19982_44348# 0.088002f
C2325 XA20.XA2.CO a_22502_43996# 0.098489f
C2326 a_12422_1390# SARN 0.014424f
C2327 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES4.B 0.430615f
C2328 XB1.TIE_L AVDD 12.9492f
C2329 XA0.CMP_OP XA5.XA1.XA4.MN1.S 0.027953f
C2330 XA1.CN0 D<1> 0.07983f
C2331 XA2.CN0 CK_SAMPLE 0.075021f
C2332 XA0.CP0 XDAC1.XC1.XRES16.B 0.028741f
C2333 XA2.XA6.MP1.S AVDD 0.092671f
C2334 XA0.CN0 VREF 0.496795f
C2335 XA6.XA6.Y XA6.XA6.MN1.S 0.026506f
C2336 XA8.XA1.XA5.MP1.S AVDD 0.087881f
C2337 XA7.XA6.Y XA7.XA6.MN3.S 0.089305f
C2338 XA5.CN0 XA5.CN1 0.050499f
C2339 XB2.XA4.GNG XDAC2.XC1.XRES8.B 0.035974f
C2340 XB1.XA4.GNG XDAC1.XC1.XRES16.B 0.098205f
C2341 a_6014_39068# AVDD 0.443169f
C2342 XA5.CP0 a_12422_45228# 0.069193f
C2343 XDAC2.XC32a<0>.XRES8.B XDAC2.XC32a<0>.XRES1A.B 0.029729f
C2344 XA0.CMP_ON a_2342_41884# 0.011704f
C2345 XA7.ENO a_17462_40124# 0.024578f
C2346 XA1.ENO a_2342_39772# 0.044989f
C2347 XA0.ENO a_3494_39772# 0.082231f
C2348 AVDD SAR_IN 0.092534f
C2349 D<2> D<1> 6.69504f
C2350 D<7> EN 0.064847f
C2351 D<4> SARN 0.034649f
C2352 D<5> VREF 1.51304f
C2353 D<6> D<8> 0.073351f
C2354 XA0.XA6.Y XA0.CP1 0.039903f
C2355 XA5.DONE AVDD 0.241164f
C2356 a_9902_40124# a_9902_39772# 0.010937f
C2357 XA3.XA2.A AVDD 2.0645f
C2358 a_11054_47692# XA4.DONE 0.023111f
C2359 a_11054_43468# VREF 0.062747f
C2360 XA6.XA8.A a_16094_47340# 0.091063f
C2361 a_2342_47692# a_2342_47340# 0.010937f
C2362 XA4.XA1.XA1.MN2.S AVDD 0.036807f
C2363 XA20.XA1.CK XA20.XA2.N1 0.331207f
C2364 XB1.TIE_L a_12422_1742# 0.157039f
C2365 XA3.CN0 XA3.CP0 3.63932f
C2366 XA2.XA1.XA1.MN2.S D<6> 0.026904f
C2367 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES8.B 0.029725f
C2368 a_n178_49100# XB1.TIE_L 0.072629f
C2369 XA4.XA11.Y XA4.XA10.Y 0.098057f
C2370 XA4.CEO XA4.XA11.MP1.S 0.010609f
C2371 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES16.B 0.05157f
C2372 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES2.B 0.033713f
C2373 XA1.ENO XA2.XA1.XA1.MP3.G 0.031841f
C2374 XA8.ENO a_21134_40828# 0.07562f
C2375 XA0.CMP_ON XA8.XA2.A 0.022245f
C2376 a_6014_43468# XA2.XA2.A 0.066256f
C2377 XDAC1.XC64a<0>.XRES1A.B SARP 3.63804f
C2378 a_22502_48220# DONE 0.071277f
C2379 XA8.XA1.XA4.LCK_N XA8.XA1.XA4.MN1.S 0.030434f
C2380 XA5.XA1.XA4.LCK_N a_13574_41180# 0.060353f
C2381 XA1.XA1.XA4.MP2.S XA1.XA1.XA4.MP1.S 0.050207f
C2382 XA0.CMP_OP a_2342_40476# 0.068716f
C2383 XA20.XA10.B XA20.XA1.CKN 0.126085f
C2384 a_n178_40476# a_n178_40124# 0.010937f
C2385 XA3.XA6.Y XA3.XA9.MN1.S 0.023798f
C2386 a_12422_45228# AVDD 0.377363f
C2387 a_23654_45404# SARN 0.02168f
C2388 a_15014_2974# a_15014_2622# 0.010937f
C2389 a_974_49452# XA0.CEO 0.040807f
C2390 a_n178_49452# XA0.XA11.Y 0.070936f
C2391 a_12422_1742# SAR_IN 0.05387f
C2392 XA3.XA1.CHL_OP XA3.CN1 0.557881f
C2393 a_11054_1390# SARN 0.032882f
C2394 a_974_48220# XA0.XA6.Y 0.066018f
C2395 a_21134_49100# AVDD 0.392086f
C2396 XDAC2.XC128a<1>.XRES1B.B SARN 3.63755f
C2397 XA0.XA1.XA4.LCK_N XA0.XA1.XA4.MN1.S 0.030434f
C2398 XA0.CMP_OP XA5.XA1.XA4.MP1.S 0.0111f
C2399 a_2342_40828# a_2342_40476# 0.010937f
C2400 XA4.XA6.MN3.S CK_SAMPLE 0.028011f
C2401 XA1.CN0 D<2> 0.079442f
C2402 XA0.CN0 SARN 0.405088f
C2403 a_7382_39420# a_7382_39068# 0.010937f
C2404 XA1.XA6.Y a_2342_46108# 0.023316f
C2405 XA6.XA6.Y XA6.CN0 0.093605f
C2406 XA4.EN XA4.ENO 0.026181f
C2407 XA5.XA1.XA5.MP1.S EN 0.03516f
C2408 a_8534_47340# a_8534_46988# 0.010937f
C2409 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES16.B 0.063821f
C2410 XDAC1.XC0.XRES8.B XDAC1.XC0.XRES2.B 0.446669f
C2411 a_12422_39420# EN 0.066018f
C2412 XA6.ENO a_18614_42588# 0.06916f
C2413 XDAC2.XC32a<0>.XRES2.B XDAC2.XC32a<0>.XRES16.B 0.470901f
C2414 XA7.XA10.Y a_18614_48572# 0.13402f
C2415 XA3.XA10.Y XA3.XA10.A 0.201839f
C2416 XA0.CMP_ON a_974_41884# 0.011248f
C2417 XA4.XA1.CHL_OP XA4.XA1.XA4.MP2.S 0.050207f
C2418 XA0.CMP_OP XA3.XA1.XA4.LCK_N 0.383512f
C2419 AVDD SAR_IP 0.092534f
C2420 D<3> D<1> 0.4436f
C2421 D<5> SARN 0.034649f
C2422 D<7> D<8> 0.073351f
C2423 D<6> VREF 1.51285f
C2424 XA4.DONE AVDD 0.241164f
C2425 XA2.XA2.A AVDD 2.06492f
C2426 a_9902_47692# XA4.DONE 0.023111f
C2427 XA3.XA8.A XA4.EN 0.144331f
C2428 XA6.XA8.A a_14942_47340# 0.127528f
C2429 XA3.XA1.XA1.MN2.S AVDD 0.036807f
C2430 XA20.XA1.CK XA20.XA3.N2 0.030618f
C2431 XA5.CN0 a_12422_46108# 0.101833f
C2432 XB1.TIE_L a_11054_1742# 0.156628f
C2433 XA4.CEO XA4.XA10.Y 0.02121f
C2434 XA1.ENO XA1.XA1.XA1.MP3.S 0.077008f
C2435 XA8.ENO a_19982_40828# 0.132757f
C2436 XA2.XA1.CHL_OP XA2.XA1.XA5.MN1.S 0.011494f
C2437 a_4862_43468# XA2.XA2.A 0.067588f
C2438 a_22502_48220# AVDD 0.391394f
C2439 XA5.XA1.XA4.LCK_N a_12422_41180# 0.023475f
C2440 XA0.CMP_OP a_974_40476# 0.067146f
C2441 XA0.CMP_ON XA6.XA1.XA1.MN2.S 0.064851f
C2442 XA4.XA1.XA1.MP3.G a_11054_40124# 0.028807f
C2443 a_6014_45228# D<6> 0.017384f
C2444 a_11054_45228# AVDD 0.377363f
C2445 XA3.XA6.Y XA3.XA8.A 0.527529f
C2446 XA8.CP0 VREF 0.610012f
C2447 XA8.XA1.XA4.MP2.S EN 0.027192f
C2448 a_n178_49452# XA0.CEO 0.023111f
C2449 XA1.ENO XA2.XA1.XA4.MN2.S 0.012065f
C2450 XA3.CP0 XA3.XA2.A 0.027978f
C2451 a_8462_686# AVDD 0.380767f
C2452 XA7.XA1.CHL_OP a_18614_44348# 0.089573f
C2453 a_n178_48220# XA0.XA6.Y 0.072725f
C2454 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES4.B 0.430615f
C2455 XDAC1.XC128b<2>.XRES1A.B SARP 3.63804f
C2456 XA0.CMP_OP XA6.XA1.XA4.MN2.S 0.025128f
C2457 a_13574_40828# XA5.XA1.XA1.MP3.G 0.066018f
C2458 XA0.XA1.XA1.MP3.G XA0.XA1.XA1.MP3.S 0.073693f
C2459 XA3.XA6.MP3.S D<5> 0.028396f
C2460 XA3.XA6.MN3.S CK_SAMPLE 0.028011f
C2461 XA1.CN0 D<3> 0.095342f
C2462 XA2.CN0 AVDD 4.36422f
C2463 XA8.XA1.XA5.MP2.S AVDD 0.033764f
C2464 a_21134_47340# XA8.ENO 0.069707f
C2465 XA5.XA1.XA4.LCK_N EN 0.038188f
C2466 XA4.CP0 a_11054_45228# 0.070763f
C2467 XA5.CN0 XA3.CN1 0.069074f
C2468 a_11054_39420# EN 0.067588f
C2469 XA7.XA10.Y a_17462_48572# 0.089492f
C2470 XA5.XA2.A XA5.XA1.XA5.MP2.S 0.050207f
C2471 XA0.CMP_ON a_n178_41884# 0.090485f
C2472 XA6.ENO a_16094_40124# 0.025674f
C2473 XA0.ENO a_974_39772# 0.054233f
C2474 D<7> VREF 1.51304f
C2475 AVDD SARP 0.164749f
C2476 D<4> D<1> 0.092293f
C2477 D<3> D<2> 6.16076f
C2478 D<6> SARN 0.034649f
C2479 XA3.DONE AVDD 0.241164f
C2480 a_8534_40124# a_8534_39772# 0.010937f
C2481 XA8.XA1.XA1.MN2.S a_19982_39772# 0.036993f
C2482 XA1.XA2.A AVDD 2.0645f
C2483 a_974_47692# a_974_47340# 0.010937f
C2484 XA3.XA6.Y XA4.EN 0.051732f
C2485 XB2.XA4.GNG XB2.XA3.B 0.379175p
C2486 XB1.M1.G a_11054_334# 0.158066f
C2487 XA1.XA1.XA1.MN2.S D<7> 0.023009f
C2488 XA3.XA1.XA1.MP2.S AVDD 0.066893f
C2489 XA8.XA11.Y a_21134_49100# 0.091063f
C2490 XA4.CEIN XA4.XA11.MP1.S 0.010771f
C2491 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES4.B 0.430615f
C2492 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES16.B 0.05157f
C2493 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES2.B 0.033713f
C2494 XA1.ENO XA1.XA1.XA1.MP3.G 0.316693f
C2495 XDAC2.XC64b<1>.XRES16.B SARN 55.2956f
C2496 a_21134_48220# AVDD 0.41338f
C2497 XA0.CMP_OP a_n178_40476# 0.09022f
C2498 XA0.CMP_ON XA5.XA1.XA1.MN2.S 0.064851f
C2499 XA8.XA1.XA1.MP3.S XA8.XA1.XA1.MP2.S 0.050207f
C2500 XA7.CP0 VREF 0.613191f
C2501 a_13862_2974# a_13862_2622# 0.010937f
C2502 XA7.ENO XA7.CN0 0.168795f
C2503 a_12422_41180# AVDD 0.39588f
C2504 a_12422_1742# SARP 0.039477f
C2505 XB1.CKN CK_SAMPLE_BSSW 0.169642f
C2506 XA7.XA1.CHL_OP a_17462_44348# 0.066439f
C2507 XA2.XA1.CHL_OP XA2.CN1 0.529833f
C2508 a_11054_1742# SAR_IP 0.05387f
C2509 XA0.CMP_OP XA5.XA1.XA4.MN2.S 0.026188f
C2510 a_974_40828# a_974_40476# 0.010937f
C2511 a_12422_40828# XA5.XA1.XA1.MP3.G 0.071498f
C2512 XA1.XA6.MN1.S CK_SAMPLE 0.053284f
C2513 XA1.XA6.MP1.S D<7> 0.016737f
C2514 XA1.CN0 D<4> 0.070487f
C2515 XA0.CN0 D<1> 0.182038f
C2516 XA0.CP1 SARP 0.334309f
C2517 a_6014_39420# a_6014_39068# 0.010937f
C2518 a_7382_47340# a_7382_46988# 0.010937f
C2519 XA6.XA1.XA5.MN2.S EN 0.016689f
C2520 XA7.XA6.Y XA7.XA6.MP3.S 0.055045f
C2521 XA8.XA1.XA4.LCK_N AVDD 0.279566f
C2522 XA2.ENO XA4.EN 1.2771f
C2523 a_19982_47340# XA8.ENO 0.067588f
C2524 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES2.B 0.033713f
C2525 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES16.B 0.05157f
C2526 XA4.CP0 a_9902_45228# 0.101124f
C2527 XA5.CN0 XA2.CN1 0.153917f
C2528 a_2342_39068# AVDD 0.442014f
C2529 XA0.ENO XA0.XA1.XA4.LCK_N 0.152052f
C2530 XA8.CEO a_23654_48220# 0.067588f
C2531 XDAC1.XC32a<0>.XRES2.B XDAC1.XC32a<0>.XRES16.B 0.470901f
C2532 XDAC1.XC32a<0>.XRES8.B XDAC1.XC32a<0>.XRES1A.B 0.029729f
C2533 AVDD EN 36.7208f
C2534 D<7> SARN 0.034649f
C2535 CK_SAMPLE VREF 2.12813f
C2536 D<4> D<2> 0.269456f
C2537 XA2.DONE AVDD 0.241164f
C2538 XA0.XA2.A AVDD 2.06497f
C2539 a_8534_47692# XA3.DONE 0.023111f
C2540 a_7382_43468# VREF 0.062747f
C2541 XA6.XA6.Y a_14942_47340# 0.011912f
C2542 XB2.CKN XB2.XA3.B 0.26479f
C2543 a_9614_1390# XB1.XA3.MP0.S 0.069705f
C2544 XA2.XA1.XA1.MP2.S AVDD 0.068123f
C2545 XA2.CN0 XA3.CP0 0.058117f
C2546 XB1.TIE_L XB1.CKN 0.066812f
C2547 XA8.XA11.Y a_19982_49100# 0.10248f
C2548 XA4.CEIN XA4.XA10.Y 0.303978f
C2549 XA3.XA11.Y XA3.XA10.Y 0.098057f
C2550 XA0.ENO XA1.XA1.XA1.MP3.G 0.126806f
C2551 XA7.ENO a_18614_40828# 0.135353f
C2552 XDAC1.XC64b<1>.XRES2.B SARP 7.01089f
C2553 XA8.CN1 XA8.XA2.A 0.703363f
C2554 a_3494_43468# XA1.XA2.A 0.066018f
C2555 XDAC2.XC64a<0>.XRES1A.B SARN 3.63804f
C2556 XA0.CMP_OP XA8.XA1.XA1.MP3.S 0.010794f
C2557 XA7.XA10.A XA7.DONE 0.045308f
C2558 XA8.XA1.XA1.MP3.G XA8.XA1.XA1.MP2.S 0.064105f
C2559 XA8.CP0 D<0> 0.177099f
C2560 XA6.CP0 VREF 0.613191f
C2561 XA3.CP0 SARP 0.046396f
C2562 XA0.CN0 XA1.CN0 6.31853f
C2563 XA7.XA1.XA4.MP1.S EN 0.027192f
C2564 XA6.ENO XA7.CN0 0.141771f
C2565 a_11054_41180# AVDD 0.39588f
C2566 a_21134_49804# a_21134_49452# 0.010937f
C2567 XA0.ENO XA1.XA1.XA4.MN2.S 0.012065f
C2568 XA2.CP0 XA2.XA2.A 0.028053f
C2569 XB2.XA4.GNG SARN 1.73183f
C2570 a_17462_49100# AVDD 0.391112f
C2571 XA6.XA1.XA5.MP2.S XA6.XA1.XA5.MP1.S 0.050207f
C2572 XA0.XA1.XA4.LCK_N XA0.XA1.XA4.MN2.S 0.030434f
C2573 XA0.CMP_OP XA4.XA1.XA4.MP1.S 0.010745f
C2574 XA0.CN0 D<2> 0.092459f
C2575 XA1.XA6.MP1.S CK_SAMPLE 0.022628f
C2576 XA0.CP1 EN 0.068864f
C2577 XA2.XA6.MP3.S D<6> 0.028396f
C2578 XA0.XA6.Y XA0.CP0 0.010942f
C2579 XA1.CN0 D<5> 0.055822f
C2580 XA5.XA1.XA5.MN2.S EN 0.016683f
C2581 XA5.CN0 XA1.CN1 0.073233f
C2582 XA4.CN0 XA4.CN1 0.050966f
C2583 XA0.CP1 XA0.XA2.A 0.03087f
C2584 XA3.CN0 XA0.CMP_ON 0.053255f
C2585 XB2.XA4.GNG XDAC2.XC1.XRES4.B 0.020556f
C2586 XB1.XA4.GNG XDAC1.XC1.XRES2.B 0.010278f
C2587 a_974_39068# AVDD 0.443169f
C2588 XA8.CEO a_22502_48220# 0.071389f
C2589 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES1A.B 0.022835f
C2590 XA4.XA1.CHL_OP XA4.XA1.XA4.MN2.S 0.062799f
C2591 XA4.XA2.A XA4.XA1.XA5.MP2.S 0.050207f
C2592 AVDD D<8> 2.0078f
C2593 D<6> D<1> 0.08931f
C2594 DONE VREF 0.089786f
C2595 D<4> D<3> 5.67288f
C2596 a_23654_47692# CK_SAMPLE 0.068482f
C2597 XA1.DONE AVDD 0.241164f
C2598 a_7382_40124# a_7382_39772# 0.010937f
C2599 XA7.XA1.XA1.MN2.S a_18614_39772# 0.036993f
C2600 a_21134_43468# AVDD 0.377891f
C2601 a_n178_47692# a_n178_47340# 0.010937f
C2602 a_7382_47692# XA3.DONE 0.023111f
C2603 a_6014_43468# VREF 0.062747f
C2604 XA2.XA8.A XA2.ENO 0.144331f
C2605 XB2.M1.G a_12422_686# 0.163985f
C2606 XB1.CKN a_9614_686# 0.114704f
C2607 XB2.CKN XB2.XA3.MP0.S 0.669708f
C2608 XA2.XA1.XA1.MN2.S AVDD 0.036807f
C2609 XA2.CN0 XA2.CP0 3.63663f
C2610 XA4.CEIN XA3.XA10.Y 0.13078f
C2611 XA3.XA11.Y XA3.XA11.MP1.S 0.054448f
C2612 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES4.B 0.430615f
C2613 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES8.B 0.477132f
C2614 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES2.B 0.015267f
C2615 XA0.ENO XA0.XA1.XA1.MP3.S 0.076247f
C2616 XA7.ENO a_17462_40828# 0.073834f
C2617 XA2.XA1.CHL_OP XA2.XA1.XA4.LCK_N 0.204048f
C2618 a_2342_43468# XA1.XA2.A 0.067827f
C2619 XDAC1.XC64a<0>.XRES16.B SARP 55.2956f
C2620 XA8.XA1.XA4.LCK_N XA8.XA1.XA4.MN2.S 0.030434f
C2621 XA0.XA1.XA4.MP2.S XA0.XA1.XA4.MP1.S 0.050207f
C2622 XA0.CMP_OP XA8.XA1.XA1.MP3.G 0.145041f
C2623 XA8.XA1.XA1.MP3.G XA8.XA1.XA1.MN2.S 0.078539f
C2624 XA3.CP0 EN 0.061409f
C2625 a_7382_45228# AVDD 0.377363f
C2626 XA5.CP0 VREF 0.613191f
C2627 XA2.CP0 SARP 0.060278f
C2628 a_15014_2974# XB2.XA2.MP0.G 0.096614f
C2629 XA0.CN0 XA0.XA6.MP1.S 0.028026f
C2630 XA5.ENO XA7.CN0 0.033243f
C2631 XB2.XA3.B AVDD 1.48564f
C2632 XA7.ENO a_19982_41884# 0.074595f
C2633 XA6.XA1.CHL_OP a_16094_44348# 0.06801f
C2634 XA1.XA1.CHL_OP XA1.CN1 0.557881f
C2635 XB1.CKN SAR_IP 0.175642f
C2636 XA20.XA10.B a_22502_48220# 0.033888f
C2637 a_16094_49100# AVDD 0.391721f
C2638 XDAC2.XC128b<2>.XRES1A.B SARN 3.63804f
C2639 XA0.CMP_OP XA4.XA1.XA4.MN1.S 0.024389f
C2640 a_n178_40828# a_n178_40476# 0.010937f
C2641 XA1.CN0 D<6> 0.06325f
C2642 XA0.CP1 D<8> 1.38522f
C2643 XA0.CN0 D<3> 0.087399f
C2644 a_4862_39420# a_4862_39068# 0.010937f
C2645 a_6014_47340# a_6014_46988# 0.010937f
C2646 XA4.XA1.XA5.MP1.S EN 0.03516f
C2647 XA7.XA1.XA5.MP1.S AVDD 0.102822f
C2648 XA6.XA1.XA4.LCK_N D<2> 0.018962f
C2649 XA1.ENO XA2.ENO 0.026181f
C2650 a_18614_47340# XA7.ENO 0.066018f
C2651 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES2.B 0.033713f
C2652 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES16.B 0.05157f
C2653 XA3.CP0 a_8534_45228# 0.102695f
C2654 XA4.CN0 XA3.CN1 0.299096f
C2655 a_7382_39420# EN 0.066018f
C2656 XA5.ENO a_14942_42588# 0.070731f
C2657 XA2.XA10.Y XA2.XA10.A 0.201839f
C2658 XDAC2.XC32a<0>.XRES8.B XDAC2.XC32a<0>.XRES16.B 0.1057f
C2659 XA0.CMP_ON XA8.XA1.XA5.MP1.S 0.025793f
C2660 XA5.ENO a_13574_40124# 0.010898f
C2661 CK_SAMPLE D<0> 0.087664f
C2662 D<6> D<2> 0.237501f
C2663 AVDD VREF 55.123604f
C2664 a_22502_47692# CK_SAMPLE 0.079928f
C2665 XA0.DONE AVDD 0.241164f
C2666 XB1.CKN a_8462_686# 0.118471f
C2667 XA1.XA1.XA1.MN2.S AVDD 0.036807f
C2668 XA4.CN0 a_11054_46108# 0.103403f
C2669 XA8.ENO XA8.XA1.CHL_OP 0.117946f
C2670 XB1.TIE_L XB2.M1.G 0.171455f
C2671 XA7.CEO a_21134_49100# 0.066018f
C2672 XA4.CEIN XA3.XA11.MP1.S 0.012048f
C2673 XA3.CN1 XA0.CMP_OP 0.273113f
C2674 XA7.CN1 XA7.XA2.A 0.703363f
C2675 XA0.ENO XA0.XA1.XA1.MP3.G 0.363295f
C2676 a_17462_48220# AVDD 0.41338f
C2677 XA0.CMP_ON XA4.XA1.XA1.MN2.S 0.064851f
C2678 XA7.XA1.XA4.LCK_N XA7.XA1.XA4.MN1.S 0.030434f
C2679 XA0.CMP_OP XA7.XA1.XA1.MP3.S 0.010682f
C2680 XA6.XA10.A XA6.DONE 0.045308f
C2681 XA2.XA9.MN1.S XA2.XA8.A 0.010335f
C2682 XA2.CP0 EN 0.06151f
C2683 a_2342_45228# D<7> 0.017384f
C2684 a_6014_45228# AVDD 0.377363f
C2685 XA3.CP0 D<8> 0.073351f
C2686 XA4.CP0 VREF 0.613191f
C2687 XA7.CP0 D<1> 0.177112f
C2688 XA1.CP0 SARP 0.177253f
C2689 a_13862_2974# XB2.XA2.MP0.G 0.067588f
C2690 XA4.ENO XA7.CN0 0.068436f
C2691 a_19982_49804# a_19982_49452# 0.010937f
C2692 XDAC2.XC64b<1>.XRES16.B XDAC2.XC64b<1>.XRES1A.B 0.467299f
C2693 XB2.XA3.MP0.S AVDD 0.183861f
C2694 XA1.CP0 XA1.XA2.A 0.027978f
C2695 XA6.XA1.CHL_OP a_14942_44348# 0.088002f
C2696 XB2.M1.G SAR_IN 0.756873f
C2697 XA6.XA1.XA4.LCK_N XA6.XA1.XA5.MN1.S 0.030434f
C2698 XA0.CMP_OP XA5.XA1.XA4.MP2.S 0.026257f
C2699 a_11054_40828# XA4.XA1.XA1.MP3.G 0.069927f
C2700 XA0.CP1 VREF 1.51285f
C2701 XA1.CN0 D<7> 0.537457f
C2702 XA0.CN0 D<4> 0.075722f
C2703 XA1.XA6.MP1.S AVDD 0.092671f
C2704 a_17462_47340# XA7.ENO 0.071277f
C2705 XA7.XA1.XA4.LCK_N AVDD 0.271288f
C2706 XA3.CP0 a_7382_45228# 0.069193f
C2707 XA4.CN0 XA2.CN1 0.668423f
C2708 a_6014_39420# EN 0.067588f
C2709 XA6.XA10.Y a_16094_48572# 0.091063f
C2710 XA3.XA1.CHL_OP XA3.XA1.XA4.MN2.S 0.062799f
C2711 XA0.CMP_ON XA8.XA1.XA5.MN1.S 0.033533f
C2712 XA5.ENO a_12422_40124# 0.024578f
C2713 D<5> D<4> 0.335782f
C2714 AVDD SARN 0.186735f
C2715 D<6> D<3> 0.088169f
C2716 CK_SAMPLE D<1> 0.106933f
C2717 a_6014_40124# a_6014_39772# 0.010937f
C2718 XA5.XA8.A a_13574_47340# 0.129098f
C2719 a_6014_47692# XA2.DONE 0.023111f
C2720 XA2.XA6.Y XA2.ENO 0.051732f
C2721 XB2.XA4.GNG a_15014_1390# 0.017291f
C2722 XA7.ENO XA8.XA1.CHL_OP 0.129613f
C2723 XA1.XA1.XA1.MP2.S AVDD 0.066893f
C2724 XA7.XA11.Y a_18614_49100# 0.104051f
C2725 XA7.CEO a_19982_49100# 0.070731f
C2726 XA2.CEO XA3.XA10.Y 0.352238f
C2727 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES2.B 0.015267f
C2728 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES8.B 0.477132f
C2729 a_974_43468# XA0.XA2.A 0.066256f
C2730 XA2.CN1 XA0.CMP_OP 0.240444f
C2731 XA6.ENO a_16094_40828# 0.075865f
C2732 XDAC2.XC64b<1>.XRES2.B SARN 7.01089f
C2733 XA1.XA1.CHL_OP XA1.XA1.XA5.MN1.S 0.011494f
C2734 a_16094_48220# AVDD 0.41338f
C2735 XA0.CMP_ON XA3.XA1.XA1.MN2.S 0.064851f
C2736 XA0.XA1.XA4.MN2.S XA0.XA1.XA4.MN1.S 0.050207f
C2737 XA0.CMP_OP XA7.XA1.XA1.MP3.G 0.142956f
C2738 XA3.XA1.XA1.MP3.G a_7382_40124# 0.028807f
C2739 XA2.XA6.Y XA2.XA8.A 0.527529f
C2740 XA1.CP0 EN 0.061409f
C2741 XA2.CP0 D<8> 0.073351f
C2742 XA3.CP0 VREF 0.629758f
C2743 XA0.CP0 SARP 0.403251f
C2744 XB1.XA2.MP0.G a_9614_2622# 0.067588f
C2745 XA6.ENO XA6.CN0 0.097278f
C2746 XA6.XA1.XA4.MP1.S EN 0.027192f
C2747 a_7382_41180# AVDD 0.39588f
C2748 XA6.ENO a_18614_41884# 0.073155f
C2749 XB2.XA3.B m3_23222_120# 0.172147f
C2750 XB1.XA3.B AVDD 1.48564f
C2751 XB1.XA4.GNG SARP 1.73183f
C2752 XA8.XA10.A a_21134_48220# 0.070424f
C2753 XA8.XA11.Y VREF 0.014797f
C2754 XA0.CMP_OP XA4.XA1.XA4.MP2.S 0.026117f
C2755 a_9902_40828# XA4.XA1.XA1.MP3.G 0.067588f
C2756 XA0.CP1 SARN 0.042322f
C2757 XA0.CN0 D<5> 0.055822f
C2758 XA1.CN0 CK_SAMPLE 0.075434f
C2759 XA3.XA6.MP3.S AVDD 0.112857f
C2760 a_3494_39420# a_3494_39068# 0.010937f
C2761 a_4862_47340# a_4862_46988# 0.010937f
C2762 XA5.XA6.Y XA5.XA6.MN1.S 0.026506f
C2763 XA6.XA6.Y XA6.XA6.MP3.S 0.055045f
C2764 XA0.ENO XA1.ENO 1.2771f
C2765 XA5.XA1.XA5.MP2.S EN 0.044153f
C2766 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES2.B 0.015267f
C2767 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES8.B 0.477132f
C2768 XA4.CN0 XA1.CN1 0.073532f
C2769 XA2.CN0 XA0.CMP_ON 0.055193f
C2770 XA4.ENO a_13574_42588# 0.06916f
C2771 a_22502_39420# AVDD 0.486332f
C2772 XA6.XA10.Y a_14942_48572# 0.13253f
C2773 XA1.XA10.Y XA1.XA10.A 0.201839f
C2774 XDAC1.XC32a<0>.XRES8.B XDAC1.XC32a<0>.XRES16.B 0.1057f
C2775 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES1A.B 0.022835f
C2776 XA0.CMP_ON XA8.XA1.XA5.MP2.S 0.010313f
C2777 XA5.CN0 XA5.XA1.XA1.MP3.G 0.016184f
C2778 CK_SAMPLE D<2> 0.106838f
C2779 D<6> D<4> 0.650867f
C2780 AVDD D<0> 1.63307f
C2781 a_21134_47692# DONE 0.047038f
C2782 a_22502_47692# AVDD 0.417082f
C2783 XA5.XA8.A a_12422_47340# 0.089492f
C2784 XA5.XA6.Y a_13574_47340# 0.011912f
C2785 a_4862_47692# XA2.DONE 0.023111f
C2786 a_17462_43468# AVDD 0.377891f
C2787 a_974_43468# D<8> 0.070763f
C2788 a_2342_43468# VREF 0.062747f
C2789 XB2.CKN a_15014_1390# 0.135393f
C2790 XA7.ENO XA7.XA1.CHL_OP 0.118011f
C2791 XA7.CN0 XA7.XA6.MP1.S 0.028026f
C2792 XA0.XA1.XA1.MP2.S AVDD 0.068123f
C2793 XA7.XA11.Y a_17462_49100# 0.089492f
C2794 XA2.XA11.Y XA2.XA11.MP1.S 0.054448f
C2795 XA2.CEO XA3.XA11.MP1.S 0.033093f
C2796 XA1.CN1 XA0.CMP_OP 0.266906f
C2797 XA6.CN1 XA6.XA2.A 0.703363f
C2798 XA6.ENO a_14942_40828# 0.132757f
C2799 a_n178_43468# XA0.XA2.A 0.067588f
C2800 XDAC1.XC64b<1>.XRES8.B SARP 27.705599f
C2801 XDAC2.XC64a<0>.XRES16.B SARN 55.2956f
C2802 XA0.CMP_OP XA6.XA1.XA1.MP3.S 0.010682f
C2803 XA0.XA6.Y a_n178_47692# 0.017683f
C2804 XA5.XA10.A XA5.DONE 0.045308f
C2805 XA7.XA1.XA1.MP3.S XA7.XA1.XA1.MP2.S 0.050207f
C2806 XA7.XA1.XA1.MP3.G XA7.XA1.XA1.MN2.S 0.078539f
C2807 XA2.XA6.Y XA2.XA9.MN1.S 0.023798f
C2808 XA6.CP0 D<2> 0.177099f
C2809 XA0.CP0 EN 0.063812f
C2810 XA1.CP0 D<8> 0.073351f
C2811 XA2.CP0 VREF 0.629107f
C2812 XA3.CP0 SARN 0.034649f
C2813 a_9614_2974# a_9614_2622# 0.010937f
C2814 XB1.XA2.MP0.G a_8462_2622# 0.072258f
C2815 a_6014_41180# AVDD 0.39588f
C2816 a_18614_49804# a_18614_49452# 0.010937f
C2817 XDAC1.XC64b<1>.XRES16.B XDAC1.XC64b<1>.XRES1A.B 0.467299f
C2818 XA0.CP0 XA0.XA2.A 0.028053f
C2819 XB2.XA3.B m3_23150_120# 0.0666f
C2820 XA5.XA1.CHL_OP a_13574_44348# 0.089573f
C2821 XA3.CN0 XA3.XA1.XA4.LCK_N 0.012456f
C2822 XB1.XA3.MP0.S AVDD 0.183861f
C2823 a_11054_1742# SARN 0.043858f
C2824 XB2.M1.G SARP 0.020328f
C2825 XA8.XA10.A a_19982_48220# 0.132671f
C2826 a_12422_49100# AVDD 0.391112f
C2827 XA8.CEO VREF 0.179573f
C2828 XDAC2.XC64a<0>.XRES1A.B XDAC2.XC1.XRES1B.B 0.62895f
C2829 XA0.CMP_OP XA3.XA1.XA4.MN1.S 0.027953f
C2830 XA0.XA6.MP1.S CK_SAMPLE 0.022425f
C2831 XA0.CN0 D<6> 0.056493f
C2832 XA2.XA6.MP3.S AVDD 0.112857f
C2833 XA5.XA6.Y XA5.XA6.MP1.S 0.055045f
C2834 a_16094_47340# XA6.ENO 0.069707f
C2835 XA4.XA1.XA5.MP2.S EN 0.044228f
C2836 XA2.CP0 a_6014_45228# 0.070763f
C2837 XB1.XA4.GNG XDAC1.XC1.XRES8.B 0.035974f
C2838 a_21134_39420# AVDD 0.472133f
C2839 XA0.CMP_ON XA8.XA1.XA4.LCK_N 0.287952f
C2840 XA0.CMP_OP XA2.XA1.XA4.LCK_N 0.375196f
C2841 XA4.ENO a_11054_40124# 0.025674f
C2842 CK_SAMPLE D<3> 0.106933f
C2843 AVDD D<1> 1.67749f
C2844 D<7> D<4> 0.013072f
C2845 D<6> D<5> 0.684738f
C2846 a_19982_47692# DONE 0.028903f
C2847 a_21134_47692# AVDD 0.393092f
C2848 a_4862_40124# a_4862_39772# 0.010937f
C2849 a_n178_43468# D<8> 0.111278f
C2850 XA0.CMP_ON EN 3.60823f
C2851 a_16094_43468# AVDD 0.377891f
C2852 a_974_43468# VREF 0.062747f
C2853 XB2.M1.G a_12422_1038# 0.16579f
C2854 XB2.CKN a_13862_1390# 0.081275f
C2855 XB1.M1.G a_11054_686# 0.163985f
C2856 XA6.ENO XA7.XA1.CHL_OP 0.13041f
C2857 XB1.TIE_L XB1.M1.G 0.170233f
C2858 XA0.XA1.XA1.MN2.S AVDD 0.036807f
C2859 XA2.XA11.Y XA2.XA10.Y 0.098057f
C2860 XA2.CEO XA2.XA11.MP1.S 0.010609f
C2861 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES8.B 0.029725f
C2862 XDAC2.X16ab.XRES16.B XDAC2.XC128b<2>.XRES16.B 0.010386f
C2863 XA1.XA1.CHL_OP XA1.XA1.XA4.LCK_N 0.204048f
C2864 XA2.XA1.CHL_OP XA2.XA1.XA5.MN2.S 0.013533f
C2865 XDAC1.XC64a<0>.XRES2.B SARP 7.01089f
C2866 XA7.XA1.XA4.LCK_N XA7.XA1.XA4.MN2.S 0.030434f
C2867 XA0.CMP_OP XA6.XA1.XA1.MP3.G 0.142977f
C2868 XA7.XA1.XA1.MP3.G XA7.XA1.XA1.MP2.S 0.064105f
C2869 XA0.CP0 D<8> 0.122159f
C2870 a_2342_45228# AVDD 0.377363f
C2871 XA1.CP0 VREF 0.629758f
C2872 XA2.CP0 SARN 0.034649f
C2873 XA7.XA1.XA4.MP2.S EN 0.027192f
C2874 XA5.XA1.CHL_OP a_12422_44348# 0.066439f
C2875 XB2.XA3.B m3_16598_280# 0.024512f
C2876 a_15014_1390# AVDD 0.380563f
C2877 a_11054_49100# AVDD 0.391721f
C2878 XA7.XA11.Y VREF 0.015777f
C2879 XA0.CMP_OP XA3.XA1.XA4.MP1.S 0.0111f
C2880 XA2.XA1.XA4.LCK_N a_4862_41884# 0.031412f
C2881 XA0.CP1 D<1> 0.094715f
C2882 XA0.XA6.MN1.S CK_SAMPLE 0.050648f
C2883 XA1.CN0 AVDD 4.4829f
C2884 a_21134_46988# D<0> 0.068712f
C2885 XA0.CN0 D<7> 0.055917f
C2886 a_2342_39420# a_2342_39068# 0.010937f
C2887 a_3494_47340# a_3494_46988# 0.010937f
C2888 a_14942_47340# XA6.ENO 0.067588f
C2889 XA5.XA1.XA4.LCK_N D<3> 0.019067f
C2890 XA4.XA1.XA4.LCK_N EN 0.038188f
C2891 XA6.XA1.XA5.MP1.S AVDD 0.102822f
C2892 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES8.B 0.477132f
C2893 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES2.B 0.015267f
C2894 XA2.CP0 a_4862_45228# 0.101124f
C2895 a_2342_39420# EN 0.066018f
C2896 XA5.XA10.Y a_13574_48572# 0.13402f
C2897 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES16.B 0.063821f
C2898 XDAC2.XC32a<0>.XRES8.B XDAC2.XC32a<0>.XRES2.B 0.446669f
C2899 XA0.CP1 XA0.XA1.XA1.MN2.S 0.026904f
C2900 XA0.CMP_ON XA7.XA1.XA5.MN1.S 0.011525f
C2901 XA3.XA1.CHL_OP XA3.XA1.XA4.MP2.S 0.050207f
C2902 XA4.XA2.A XA4.XA1.XA5.MN2.S 0.050207f
C2903 CK_SAMPLE D<4> 0.106838f
C2904 AVDD D<2> 1.67477f
C2905 D<7> D<5> 0.290865f
C2906 XA1.XA8.A XA1.ENO 0.144331f
C2907 XA20.XA10.A XA20.XA1.CKN 0.321724f
C2908 a_3494_47692# XA1.DONE 0.023111f
C2909 XA0.CMP_ON D<8> 0.180502f
C2910 XA6.ENO XA6.XA1.CHL_OP 0.117946f
C2911 XA20.XA1.MP0.S AVDD 0.428745f
C2912 XA6.CEO a_18614_49100# 0.0733f
C2913 XA2.CEO XA2.XA10.Y 0.02121f
C2914 XA5.CN1 XA5.XA2.A 0.703363f
C2915 XA5.ENO a_13574_40828# 0.135353f
C2916 a_12422_48220# AVDD 0.41338f
C2917 XA8.XA10.A VREF 0.015558f
C2918 XA4.XA1.XA4.LCK_N a_11054_41180# 0.023475f
C2919 XA0.CMP_ON XA2.XA1.XA1.MN2.S 0.064851f
C2920 XA0.CMP_OP XA5.XA1.XA1.MP3.S 0.010682f
C2921 XA20.XA10.B a_23654_47692# 0.066264f
C2922 XA4.XA10.A XA4.DONE 0.045308f
C2923 XA2.XA1.XA1.MP3.G a_6014_40124# 0.028807f
C2924 XA0.CP0 VREF 0.629107f
C2925 XA5.CP0 D<3> 0.177112f
C2926 XA3.CP0 D<1> 0.011917f
C2927 a_974_45228# AVDD 0.377363f
C2928 XA1.CP0 SARN 0.034649f
C2929 a_8462_2974# a_8462_2622# 0.010937f
C2930 a_15014_3326# a_15014_2974# 0.010937f
C2931 XA6.XA1.XA4.MP2.S EN 0.027192f
C2932 a_17462_49804# a_17462_49452# 0.010937f
C2933 XDAC2.XC64b<1>.XRES2.B XDAC2.XC64b<1>.XRES1A.B 0.015267f
C2934 XB1.M1.G SAR_IP 0.755165f
C2935 XB2.XA3.B m3_16526_280# 0.024512f
C2936 XA7.XA10.A a_18614_48220# 0.134161f
C2937 XA7.CEO VREF 0.019575f
C2938 XDAC1.XC64a<0>.XRES1A.B XDAC1.XC1.XRES1B.B 0.62895f
C2939 XA6.XA1.XA5.MN2.S XA6.XA1.XA5.MN1.S 0.050207f
C2940 XA0.CMP_OP XA4.XA1.XA4.MN2.S 0.025128f
C2941 a_8534_40828# XA3.XA1.XA1.MP3.G 0.066018f
C2942 XA0.XA6.MP1.S AVDD 0.092671f
C2943 XA0.CN0 CK_SAMPLE 0.075021f
C2944 a_974_39420# EN 0.067588f
C2945 XA5.XA10.Y a_12422_48572# 0.089492f
C2946 CK_SAMPLE D<5> 0.106933f
C2947 AVDD D<3> 1.67749f
C2948 D<7> D<6> 1.44168f
C2949 XA1.CN0 XDAC2.XC64a<0>.XRES16.B 0.025998f
C2950 a_3494_40124# a_3494_39772# 0.010937f
C2951 XA6.XA1.XA1.MN2.S a_14942_39772# 0.036993f
C2952 XA1.XA6.Y XA1.ENO 0.051732f
C2953 XA4.XA8.A a_11054_47340# 0.091063f
C2954 a_2342_47692# XA1.DONE 0.023111f
C2955 XA0.CMP_ON VREF 0.116975f
C2956 XB1.CKN XB1.XA3.B 0.26479f
C2957 XB2.M1.G XB2.XA3.B 0.016334f
C2958 XA5.ENO XA6.XA1.CHL_OP 0.129613f
C2959 XA1.CN0 XA3.CP0 0.058178f
C2960 XA0.CP1 a_974_45228# 0.017384f
C2961 a_21134_40476# AVDD 0.362621f
C2962 XA6.XA11.Y a_16094_49100# 0.091063f
C2963 XA6.CEO a_17462_49100# 0.07472f
C2964 XA1.CEO XA2.XA11.MP1.S 0.010771f
C2965 XDAC2.XC128b<2>.XRES1A.B XDAC2.XC128a<1>.XRES1B.B 0.62895f
C2966 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES8.B 0.029725f
C2967 XDAC1.X16ab.XRES16.B XDAC1.XC128b<2>.XRES16.B 0.010386f
C2968 XA5.ENO a_12422_40828# 0.073834f
C2969 XA1.XA1.CHL_OP XA1.XA1.XA5.MN2.S 0.013533f
C2970 XDAC2.XC64b<1>.XRES8.B SARN 27.705599f
C2971 a_11054_48220# AVDD 0.41338f
C2972 XA7.XA10.A VREF 0.015839f
C2973 XA4.XA1.XA4.LCK_N a_9902_41180# 0.060353f
C2974 XA0.CMP_ON XA1.XA1.XA1.MN2.S 0.064851f
C2975 XA0.CMP_OP XA5.XA1.XA1.MP3.G 0.142956f
C2976 XA20.XA10.B a_22502_47692# 0.100549f
C2977 XA6.XA1.XA1.MP3.S XA6.XA1.XA1.MP2.S 0.050207f
C2978 a_21134_46108# VREF 0.031902f
C2979 XA3.CP0 D<2> 0.016387f
C2980 XA0.CP0 SARN 0.034649f
C2981 XA0.CP1 XA0.XA6.MP1.S 0.016737f
C2982 a_2342_41180# AVDD 0.39588f
C2983 XA4.XA1.CHL_OP a_11054_44348# 0.06801f
C2984 XA5.ENO a_14942_41884# 0.074595f
C2985 XB1.M1.G SARP 0.308182f
C2986 XB2.XA3.B m3_23222_1080# 0.172147f
C2987 XA6.XA11.Y VREF 0.015286f
C2988 XA0.XA10.A XA0.XA9.MN1.S 0.073313f
C2989 XA7.XA10.A a_17462_48220# 0.068853f
C2990 XA0.CMP_OP XA3.XA1.XA4.MN2.S 0.026188f
C2991 XA20.XA2.N1 a_22502_40828# 0.023111f
C2992 a_7382_40828# XA3.XA1.XA1.MP3.G 0.071498f
C2993 XA2.XA6.MN3.S CK_SAMPLE 0.028011f
C2994 a_974_39420# a_974_39068# 0.010937f
C2995 a_2342_47340# a_2342_46988# 0.010937f
C2996 XA5.XA6.Y XA5.CN0 0.093605f
C2997 a_13574_47340# XA5.ENO 0.066018f
C2998 XA3.XA1.XA5.MP1.S EN 0.03516f
C2999 XA7.XA1.XA5.MP2.S AVDD 0.038567f
C3000 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES8.B 0.029725f
C3001 XA1.CP0 a_3494_45228# 0.102695f
C3002 XA4.EN a_9902_42588# 0.070731f
C3003 a_n178_39420# EN 0.071606f
C3004 a_17462_39420# AVDD 0.470715f
C3005 XA0.XA10.Y XA0.XA10.A 0.201839f
C3006 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES16.B 0.063821f
C3007 XDAC1.XC32a<0>.XRES8.B XDAC1.XC32a<0>.XRES2.B 0.446669f
C3008 XA0.CMP_ON XA7.XA1.XA4.LCK_N 0.284482f
C3009 XA2.XA1.CHL_OP XA2.XA1.XA4.MP2.S 0.050207f
C3010 XA0.CMP_OP XA1.XA1.XA4.LCK_N 0.383512f
C3011 XA3.XA2.A XA3.XA1.XA5.MN2.S 0.050207f
C3012 XA4.EN a_8534_40124# 0.010898f
C3013 CK_SAMPLE D<6> 0.106838f
C3014 AVDD D<4> 1.67477f
C3015 a_17462_47692# AVDD 0.395235f
C3016 XA4.XA8.A a_9902_47340# 0.127528f
C3017 XA8.CN1 EN 0.024032f
C3018 a_12422_43468# AVDD 0.377891f
C3019 a_12422_1742# a_12422_1390# 0.010937f
C3020 XB1.CKN XB1.XA3.MP0.S 0.669708f
C3021 XB1.XA4.GNG XB1.XA3.B 0.379175p
C3022 XA1.CN0 XA2.CP0 0.064892f
C3023 XA5.ENO XA5.XA1.CHL_OP 0.118011f
C3024 XA20.XA1.CK XA20.XA2.VMR 0.380687f
C3025 XB1.TIE_L XB2.XA1.Y 0.047823f
C3026 XA6.XA11.Y a_14942_49100# 0.10248f
C3027 XA6.CEO a_16094_49100# 0.015625f
C3028 XA1.CEO XA2.XA10.Y 0.303978f
C3029 XA1.XA11.Y XA1.XA10.Y 0.098057f
C3030 XA4.CN1 XA4.XA2.A 0.703363f
C3031 XA8.XA1.CHL_OP a_19982_42588# 0.01727f
C3032 XDAC1.XC64b<1>.XRES4.B SARP 13.9307f
C3033 XDAC1.XC64b<1>.XRES16.B D<7> 0.027052f
C3034 XA6.XA10.A VREF 0.015839f
C3035 XDAC2.XC64a<0>.XRES2.B SARN 7.01089f
C3036 XA0.CMP_OP XA4.XA1.XA1.MP3.S 0.010682f
C3037 XA3.XA10.A XA3.DONE 0.045308f
C3038 XA6.XA1.XA1.MP3.G XA6.XA1.XA1.MP2.S 0.064105f
C3039 XA1.XA8.A XA1.XA9.MN1.S 0.010335f
C3040 XA1.XA6.Y XA2.XA6.Y 0.046858f
C3041 XA3.CP0 D<3> 0.026145f
C3042 XA4.CP0 D<4> 0.177099f
C3043 XA8.CP0 CK_SAMPLE 0.038932f
C3044 XA1.CP0 D<1> 0.087788f
C3045 a_13862_3326# a_13862_2974# 0.010937f
C3046 XA5.XA1.XA4.MP1.S EN 0.027192f
C3047 a_974_41180# AVDD 0.39588f
C3048 a_16094_49804# a_16094_49452# 0.010937f
C3049 XDAC1.XC64b<1>.XRES2.B XDAC1.XC64b<1>.XRES1A.B 0.015267f
C3050 XA4.XA1.CHL_OP a_9902_44348# 0.088002f
C3051 XB2.XA1.Y SAR_IN 0.023477f
C3052 XB2.M1.G SARN 0.410932f
C3053 XB2.XA3.B m3_23150_1080# 0.0666f
C3054 a_7382_49100# AVDD 0.391112f
C3055 XA6.CEO VREF 0.367402f
C3056 XA0.XA10.A XA0.XA6.Y 0.205884f
C3057 XA0.CMP_OP XA2.XA1.XA4.MP1.S 0.010745f
C3058 XA0.CN0 AVDD 4.3574f
C3059 XA1.XA6.MP3.S D<7> 0.028396f
C3060 XA1.XA6.MN3.S CK_SAMPLE 0.028011f
C3061 XA6.XA6.Y XA6.XA6.MN3.S 0.089305f
C3062 a_12422_47340# XA5.ENO 0.071277f
C3063 XA3.XA1.XA4.LCK_N EN 0.038188f
C3064 XA6.XA1.XA5.MP2.S AVDD 0.038567f
C3065 XA1.CP0 a_2342_45228# 0.069193f
C3066 XA3.CN0 XA3.CN1 3.1969f
C3067 XA20.XA1.CK XA0.CMP_OP 0.045599f
C3068 XB1.XA4.GNG XDAC1.XC1.XRES4.B 0.020556f
C3069 a_21134_39772# EN 0.071657f
C3070 a_16094_39420# AVDD 0.471851f
C3071 XA4.EN a_7382_40124# 0.024578f
C3072 XA4.CN0 XA4.XA1.XA1.MP3.G 0.021257f
C3073 CK_SAMPLE D<7> 0.106933f
C3074 AVDD D<5> 1.5988f
C3075 XA8.XA1.XA4.MP2.S XA8.XA1.XA4.MP1.S 0.050207f
C3076 a_16094_47692# AVDD 0.395235f
C3077 XA5.XA1.XA1.MN2.S a_13574_39772# 0.036993f
C3078 a_2342_40124# a_2342_39772# 0.010937f
C3079 XA0.XA8.A XA0.ENO 0.144331f
C3080 a_974_47692# XA0.DONE 0.023111f
C3081 XA7.CN1 EN 0.024032f
C3082 a_11054_43468# AVDD 0.377891f
C3083 XB1.M1.G a_11054_1038# 0.16579f
C3084 XA1.CN0 XA1.CP0 3.78756f
C3085 XA4.ENO XA5.XA1.CHL_OP 0.13041f
C3086 XA20.XA1.CK XA20.XA2.CO 0.530644f
C3087 XB1.TIE_L a_12422_2094# 0.157781f
C3088 XA1.CEO XA1.XA10.Y 0.13078f
C3089 XA1.XA11.Y XA1.XA11.MP1.S 0.054448f
C3090 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES4.B 0.430615f
C3091 XDAC1.XC128b<2>.XRES1A.B XDAC1.XC128a<1>.XRES1B.B 0.62895f
C3092 XA8.CN1 a_21134_43468# 0.070763f
C3093 XA4.ENO a_11054_40828# 0.075865f
C3094 XA5.XA10.A VREF 0.015839f
C3095 XDAC1.XC64a<0>.XRES8.B SARP 27.705599f
C3096 XA0.CMP_OP XA4.XA1.XA1.MP3.G 0.142977f
C3097 XA6.XA1.XA1.MP3.G XA6.XA1.XA1.MN2.S 0.078539f
C3098 XA1.XA6.Y XA1.XA9.MN1.S 0.023798f
C3099 XA0.CP0 D<1> 0.099397f
C3100 XA1.CP0 D<2> 0.086501f
C3101 a_21134_46108# D<0> 0.011483f
C3102 XA3.CP0 D<4> 3.05097f
C3103 XA7.CP0 CK_SAMPLE 0.054325f
C3104 a_22502_45404# AVDD 0.416863f
C3105 XA0.CP1 XA0.CN0 0.475911f
C3106 XA4.ENO a_13574_41884# 0.073155f
C3107 a_12422_2094# SAR_IN 0.05378f
C3108 XB2.XA3.B m3_16598_1240# 0.024512f
C3109 a_6014_49100# AVDD 0.391721f
C3110 XA5.XA11.Y VREF 0.015777f
C3111 XA6.XA10.A a_16094_48220# 0.070424f
C3112 XA5.XA1.XA4.LCK_N XA5.XA1.XA5.MN1.S 0.030434f
C3113 XA6.XA1.XA5.MN2.S XA6.XA1.XA4.LCK_N 0.010898f
C3114 XA1.XA1.XA4.LCK_N a_3494_41884# 0.031412f
C3115 XA0.CMP_OP XA2.XA1.XA4.MN1.S 0.024389f
C3116 a_17462_46988# D<1> 0.070283f
C3117 XA0.CP1 D<5> 0.792851f
C3118 a_n178_39420# a_n178_39068# 0.010937f
C3119 a_974_47340# a_974_46988# 0.010937f
C3120 XA4.XA1.XA5.MN2.S EN 0.016689f
C3121 XA6.XA1.XA4.LCK_N AVDD 0.271451f
C3122 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES8.B 0.029725f
C3123 XA3.CN0 XA2.CN1 0.152577f
C3124 XA2.ENO a_8534_42588# 0.06916f
C3125 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES16.B 0.05157f
C3126 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES2.B 0.033713f
C3127 XA20.XA2.N1 XA20.XA2.N2 0.474658f
C3128 AVDD D<6> 1.59889f
C3129 a_n178_47692# XA0.DONE 0.023111f
C3130 XA4.XA6.Y a_9902_47340# 0.011912f
C3131 XA7.XA8.A XA7.DONE 0.1303f
C3132 XA0.CMP_ON D<1> 0.064523f
C3133 XA6.CN1 EN 0.024032f
C3134 XA8.CN1 VREF 0.614849f
C3135 XB2.CKN XB2.XA4.GNG 0.142777f
C3136 a_11054_1742# a_11054_1390# 0.010937f
C3137 XA4.ENO XA4.XA1.CHL_OP 0.117946f
C3138 XB1.TIE_L a_11054_2094# 0.15737f
C3139 XA0.CN0 XA3.CP0 0.127416f
C3140 a_17462_40476# AVDD 0.362093f
C3141 XA5.CEO a_16094_49100# 0.066018f
C3142 XA1.CEO XA1.XA11.MP1.S 0.012048f
C3143 XA3.CN1 XA3.XA2.A 0.749811f
C3144 XA8.CN1 a_19982_43468# 0.107905f
C3145 XA7.XA1.CHL_OP a_18614_42588# 0.01727f
C3146 XA4.ENO a_9902_40828# 0.132757f
C3147 XA0.XA1.CHL_OP XA0.XA1.XA5.MN1.S 0.011494f
C3148 a_7382_48220# AVDD 0.41338f
C3149 XA4.XA10.A VREF 0.015839f
C3150 XA0.CMP_ON XA0.XA1.XA1.MN2.S 0.064851f
C3151 XA0.CMP_OP XA3.XA1.XA1.MP3.S 0.010682f
C3152 XA2.XA10.A XA2.DONE 0.045308f
C3153 a_22502_48220# XA20.XA10.A 0.023111f
C3154 a_17462_46108# VREF 0.031953f
C3155 XA1.CP0 D<3> 0.086573f
C3156 XA0.CP0 D<2> 0.098065f
C3157 XA2.CP0 D<4> 0.224159f
C3158 XA1.XA6.Y XA1.XA8.A 0.527529f
C3159 XA3.CP0 D<5> 6.69167f
C3160 XA6.CP0 CK_SAMPLE 0.054172f
C3161 XA8.CP0 AVDD 2.11017f
C3162 XA8.XA1.XA4.MP1.S AVDD 0.091926f
C3163 a_14942_49804# a_14942_49452# 0.010937f
C3164 XDAC2.XC64b<1>.XRES8.B XDAC2.XC64b<1>.XRES1A.B 0.029729f
C3165 XDAC2.XC64b<1>.XRES2.B XDAC2.XC64b<1>.XRES16.B 0.470901f
C3166 XA3.XA1.CHL_OP a_8534_44348# 0.089573f
C3167 XB2.XA3.B m3_16526_1240# 0.024512f
C3168 a_8462_1390# AVDD 0.380563f
C3169 XA5.CEO VREF 0.018904f
C3170 a_23654_48572# a_23654_48220# 0.010937f
C3171 XA6.XA10.A a_14942_48220# 0.132671f
C3172 XA0.CMP_OP XA3.XA1.XA4.MP2.S 0.026257f
C3173 a_6014_40828# XA2.XA1.XA1.MP3.G 0.069927f
C3174 XA0.CP1 D<6> 0.134808f
C3175 a_11054_47340# XA4.ENO 0.069707f
C3176 XA3.XA1.XA5.MN2.S EN 0.016683f
C3177 XA1.CN0 XA0.CMP_ON 0.053255f
C3178 XA3.CN0 XA1.CN1 0.077513f
C3179 XA0.CP0 a_974_45228# 0.070763f
C3180 XA4.XA10.Y a_11054_48572# 0.091063f
C3181 XA2.XA1.CHL_OP XA2.XA1.XA4.MN2.S 0.062799f
C3182 XA3.XA2.A XA3.XA1.XA5.MP2.S 0.050207f
C3183 XA2.ENO a_6014_40124# 0.025674f
C3184 XA8.ENO XA8.XA1.XA1.MP2.S 0.150467f
C3185 AVDD D<7> 1.5988f
C3186 DONE CK_SAMPLE 0.399423f
C3187 a_974_40124# a_974_39772# 0.010937f
C3188 XA5.CN1 EN 0.024032f
C3189 XA0.CMP_ON D<2> 0.06424f
C3190 XA7.XA6.Y XA7.DONE 0.014904f
C3191 XA7.CN1 VREF 0.618029f
C3192 XB2.M1.G a_15014_1390# 0.034677f
C3193 XA4.EN XA4.XA1.CHL_OP 0.129613f
C3194 XA8.ENO XA20.XA2.VMR 0.159182f
C3195 XA6.CN0 XA7.CN0 7.16663f
C3196 XA0.CN0 XA2.CP0 0.058178f
C3197 a_16094_40476# AVDD 0.362177f
C3198 XA0.CEO XA1.XA10.Y 0.352238f
C3199 XA5.CEO a_14942_49100# 0.070731f
C3200 XA5.XA11.Y a_13574_49100# 0.104051f
C3201 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES4.B 0.430615f
C3202 XDAC2.XC64b<1>.XRES4.B SARN 13.9307f
C3203 a_6014_48220# AVDD 0.41338f
C3204 XA3.XA10.A VREF 0.015839f
C3205 XA3.XA1.XA4.LCK_N a_8534_41180# 0.060353f
C3206 XA0.CMP_OP XA3.XA1.XA1.MP3.G 0.142956f
C3207 XA1.XA1.XA1.MP3.G a_2342_40124# 0.028807f
C3208 a_16094_46108# VREF 0.031953f
C3209 XA0.CP0 D<3> 0.098764f
C3210 XA1.CP0 D<4> 0.118392f
C3211 XA2.CP0 D<5> 3.80406f
C3212 XA5.CP0 CK_SAMPLE 0.054325f
C3213 XA7.CP0 AVDD 2.04538f
C3214 XA3.CP0 D<6> 0.084511f
C3215 XA5.ENO XA5.CN0 0.168549f
C3216 XA4.XA1.XA4.MP1.S EN 0.027192f
C3217 XA3.XA1.CHL_OP a_7382_44348# 0.066439f
C3218 XB1.M1.G SARN 0.175565f
C3219 XDAC2.XC128b<2>.XRES16.B XDAC2.XC128a<1>.XRES16.B 0.010386f
C3220 XB2.XA3.B m3_23222_2040# 0.172147f
C3221 XB2.XA4.GNG AVDD 2.51656f
C3222 a_11054_2094# SAR_IP 0.05378f
C3223 a_12422_2094# SARP 0.041929f
C3224 XA4.XA11.Y VREF 0.015286f
C3225 XA5.XA1.XA5.MN2.S XA5.XA1.XA5.MN1.S 0.050207f
C3226 XA0.CMP_OP XA2.XA1.XA4.MP2.S 0.026117f
C3227 a_4862_40828# XA2.XA1.XA1.MP3.G 0.067588f
C3228 XA0.CP1 D<7> 0.792962f
C3229 XA1.XA6.MP3.S AVDD 0.112857f
C3230 a_16094_46988# D<2> 0.068712f
C3231 XA0.XA6.MN3.S CK_SAMPLE 0.028011f
C3232 XA2.XA1.XA5.MP1.S EN 0.03516f
C3233 a_n178_47340# a_n178_46988# 0.010937f
C3234 XA4.XA6.Y XA4.XA6.MP1.S 0.055045f
C3235 a_9902_47340# XA4.ENO 0.067588f
C3236 XA5.XA1.XA5.MP1.S AVDD 0.102822f
C3237 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES4.B 0.430615f
C3238 XA8.ENO XA0.CMP_OP 0.359924f
C3239 XA2.CN0 XA3.CN1 3.54207f
C3240 XA20.XA4.MP0.S XA20.XA2.VMR 0.095491f
C3241 XA0.CP0 a_n178_45228# 0.101124f
C3242 a_17462_39772# EN 0.073293f
C3243 a_12422_39420# AVDD 0.470715f
C3244 XA4.XA10.Y a_9902_48572# 0.13253f
C3245 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES16.B 0.05157f
C3246 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES2.B 0.033713f
C3247 XA0.CMP_ON XA6.XA1.XA5.MN1.S 0.011062f
C3248 XA8.ENO XA8.XA1.XA1.MN2.S 0.040111f
C3249 AVDD CK_SAMPLE 5.08392f
C3250 a_12422_47692# AVDD 0.395235f
C3251 XA8.XA8.A VREF 0.027267f
C3252 XA8.CN1 D<0> 0.590469f
C3253 XA4.CN1 EN 0.024032f
C3254 XA0.CMP_ON D<3> 0.064471f
C3255 XA6.CN1 VREF 0.618029f
C3256 a_7382_43468# AVDD 0.377891f
C3257 XA3.CN1 SARP 0.06043f
C3258 XB2.XA4.MN1.S XB2.CKN 0.011708f
C3259 XB1.M1.G XB1.XA3.B 0.016334f
C3260 XA8.ENO XA20.XA2.CO 0.012697f
C3261 XA4.EN XA3.XA1.CHL_OP 0.118011f
C3262 XA6.CN0 XA6.XA6.MP1.S 0.028026f
C3263 XA3.CN0 a_7382_46108# 0.101833f
C3264 XA0.CN0 XA1.CP0 0.112241f
C3265 XA8.XA1.XA1.MP3.G EN 0.145323f
C3266 XA0.CEO XA1.XA11.MP1.S 0.033093f
C3267 XA0.XA11.Y XA0.XA11.MP1.S 0.054448f
C3268 XA5.XA11.Y a_12422_49100# 0.089492f
C3269 XA2.CN1 XA2.XA2.A 0.748414f
C3270 XA7.CN1 a_18614_43468# 0.109463f
C3271 XA4.EN a_8534_40828# 0.135353f
C3272 XDAC1.XC64b<1>.XRES1B.B SARP 3.63755f
C3273 XA2.XA10.A VREF 0.015839f
C3274 XDAC2.XC64a<0>.XRES8.B SARN 27.705599f
C3275 XA3.XA1.XA4.LCK_N a_7382_41180# 0.023475f
C3276 XA0.CMP_OP XA2.XA1.XA1.MP3.S 0.010682f
C3277 XA1.XA10.A XA1.DONE 0.045308f
C3278 a_21134_48220# XA8.XA6.Y 0.066018f
C3279 XA5.XA1.XA1.MP3.S XA5.XA1.XA1.MP2.S 0.050207f
C3280 XA5.XA1.XA1.MP3.G XA5.XA1.XA1.MN2.S 0.078539f
C3281 XA6.CP0 AVDD 2.04562f
C3282 XA1.CP0 D<5> 0.483256f
C3283 XA0.CP0 D<4> 0.109242f
C3284 XA4.CP0 CK_SAMPLE 0.054172f
C3285 XA2.CP0 D<6> 7.01117f
C3286 XA4.ENO XA5.CN0 0.064699f
C3287 XA8.XA1.XA4.MP2.S AVDD 0.046398f
C3288 a_13574_49804# a_13574_49452# 0.010937f
C3289 XDAC1.XC64b<1>.XRES2.B XDAC1.XC64b<1>.XRES16.B 0.470901f
C3290 XDAC1.XC64b<1>.XRES8.B XDAC1.XC64b<1>.XRES1A.B 0.029729f
C3291 XA20.XA3.N2 XA20.XA2.N1 0.440586f
C3292 XB2.XA3.B m3_23150_2040# 0.0666f
C3293 XB2.CKN AVDD 2.35133f
C3294 a_2342_49100# AVDD 0.391112f
C3295 XA4.CEO VREF 0.367402f
C3296 a_22502_48572# a_22502_48220# 0.010937f
C3297 XA5.XA10.A a_13574_48220# 0.134161f
C3298 XDAC2.XC64a<0>.XRES16.B XDAC2.XC64a<0>.XRES1A.B 0.467299f
C3299 XA0.CMP_OP XA1.XA1.XA4.MN1.S 0.027953f
C3300 XA0.XA6.MP3.S AVDD 0.112857f
C3301 XA0.CP1 CK_SAMPLE 0.106828f
C3302 XA4.XA6.Y XA4.XA6.MN1.S 0.026506f
C3303 XA5.XA6.Y XA5.XA6.MN3.S 0.089305f
C3304 XA5.XA1.XA4.LCK_N AVDD 0.271288f
C3305 XA7.CN0 XA7.XA1.CHL_OP 0.037394f
C3306 XA7.ENO XA0.CMP_OP 0.819174f
C3307 XA2.CN0 XA2.CN1 3.16895f
C3308 a_16094_39772# EN 0.071722f
C3309 a_11054_39420# AVDD 0.471851f
C3310 XA7.ENO XA8.XA1.XA1.MN2.S 0.030034f
C3311 XA2.XA2.A XA2.XA1.XA5.MP2.S 0.050207f
C3312 XA1.XA1.CHL_OP XA1.XA1.XA4.MN2.S 0.062799f
C3313 XA8.XA1.CHL_OP a_21134_41884# 0.023777f
C3314 AVDD DONE 1.55845f
C3315 XA8.XA1.XA4.MN2.S XA8.XA1.XA4.MN1.S 0.050207f
C3316 a_11054_47692# AVDD 0.395235f
C3317 a_n178_40124# a_n178_39772# 0.010937f
C3318 XA3.CN1 EN 0.09808f
C3319 XA0.CMP_ON D<4> 0.064267f
C3320 XA6.XA8.A XA6.DONE 0.1303f
C3321 XA3.XA8.A a_8534_47340# 0.129098f
C3322 XA5.CN1 VREF 0.618029f
C3323 a_6014_43468# AVDD 0.377891f
C3324 XA2.CN1 SARP 0.050102f
C3325 XB1.CKN a_9614_1390# 0.082845f
C3326 XB2.M1.G a_12422_1390# 0.070815f
C3327 XA2.ENO XA3.XA1.CHL_OP 0.13041f
C3328 XA0.CN0 XA0.CP0 6.35579f
C3329 XA0.CEO XA0.XA11.MP1.S 0.010609f
C3330 XA0.XA11.Y XA0.XA10.Y 0.098057f
C3331 XA0.XA1.CHL_OP XA0.XA1.XA4.LCK_N 0.204048f
C3332 XA7.CN1 a_17462_43468# 0.069193f
C3333 XA4.EN a_7382_40828# 0.073834f
C3334 XA1.XA10.A VREF 0.015839f
C3335 XDAC1.XC64a<0>.XRES4.B SARP 13.9307f
C3336 XA0.CMP_OP XA2.XA1.XA1.MP3.G 0.142977f
C3337 a_19982_48220# XA8.XA6.Y 0.072725f
C3338 XA5.XA1.XA1.MP3.G XA5.XA1.XA1.MP2.S 0.064105f
C3339 XA5.CP0 AVDD 2.04538f
C3340 a_17462_46108# D<1> 0.011483f
C3341 XA0.CP0 D<5> 0.601791f
C3342 XA2.CP0 D<7> 1.26437f
C3343 XA1.CP0 D<6> 6.33012f
C3344 XA3.CP0 CK_SAMPLE 0.054325f
C3345 a_9614_2974# XB1.XA2.MP0.G 0.066018f
C3346 XA0.CP1 XA0.XA6.MP3.S 0.028396f
C3347 XA5.XA1.XA4.MP2.S EN 0.027192f
C3348 XA2.XA1.CHL_OP a_6014_44348# 0.06801f
C3349 XA4.EN a_9902_41884# 0.074595f
C3350 XDAC1.XC128b<2>.XRES16.B XDAC1.XC128a<1>.XRES16.B 0.010386f
C3351 XB2.XA4.GNG m3_23222_120# 0.049023f
C3352 XB2.XA3.B m3_16598_2200# 0.024512f
C3353 a_974_49100# AVDD 0.391721f
C3354 XA3.XA11.Y VREF 0.015777f
C3355 XA5.XA10.A a_12422_48220# 0.068853f
C3356 XA5.XA1.XA5.MN2.S XA5.XA1.XA4.LCK_N 0.010898f
C3357 XA0.CMP_OP XA1.XA1.XA4.MP1.S 0.0111f
C3358 a_21134_39772# a_21134_39420# 0.010937f
C3359 XA4.XA1.XA4.LCK_N D<4> 0.018962f
C3360 XA4.XA6.Y XA4.CN0 0.093605f
C3361 XA3.XA1.XA5.MP2.S EN 0.044153f
C3362 a_8534_47340# XA4.EN 0.066018f
C3363 XA20.XA1.CKN XA20.XA1.CK 1.59187f
C3364 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES4.B 0.430615f
C3365 XA1.ENO a_4862_42588# 0.070731f
C3366 XA6.ENO XA0.CMP_OP 0.6934f
C3367 XA2.CN0 XA1.CN1 0.083981f
C3368 XA0.CN0 XA0.CMP_ON 0.055193f
C3369 XA3.XA10.Y a_8534_48572# 0.13402f
C3370 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES8.B 0.477132f
C3371 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES2.B 0.015267f
C3372 XA7.ENO XA7.XA1.XA1.MN2.S 0.104122f
C3373 XA1.ENO a_3494_40124# 0.010898f
C3374 XA8.XA1.CHL_OP a_19982_41884# 0.040867f
C3375 XA0.XA6.Y a_974_46988# 0.023982f
C3376 XA2.CN1 EN 0.099922f
C3377 XA0.CMP_ON D<5> 0.056276f
C3378 XA3.CN1 D<8> 1.71572f
C3379 XA3.XA6.Y a_8534_47340# 0.011912f
C3380 XA3.XA8.A a_7382_47340# 0.089492f
C3381 XA4.CN1 VREF 0.618029f
C3382 XA7.CN1 D<1> 0.62381f
C3383 XA1.CN1 SARP 0.042583f
C3384 XB1.CKN a_8462_1390# 0.135393f
C3385 XA2.ENO XA2.XA1.CHL_OP 0.117946f
C3386 a_12422_40476# AVDD 0.362093f
C3387 XA7.XA1.XA1.MP3.G EN 0.145483f
C3388 XA0.CEO XA0.XA10.Y 0.02121f
C3389 XA0.XA11.Y XB1.TIE_L 0.222689f
C3390 XA4.CEO a_13574_49100# 0.0733f
C3391 XA0.XA1.CHL_OP XA0.XA1.XA5.MN2.S 0.013533f
C3392 XA1.CN1 XA1.XA2.A 0.749811f
C3393 XA6.XA1.CHL_OP a_14942_42588# 0.01727f
C3394 a_2342_48220# AVDD 0.41338f
C3395 XA0.XA10.A VREF 0.015839f
C3396 XA6.XA1.XA4.LCK_N XA6.XA1.XA4.MN1.S 0.030434f
C3397 XA0.CMP_OP XA1.XA1.XA1.MP3.S 0.010682f
C3398 XA0.XA10.A XA0.DONE 0.045308f
C3399 XA0.XA1.XA1.MP3.G a_974_40124# 0.028807f
C3400 XA4.CP0 AVDD 2.04562f
C3401 a_12422_46108# VREF 0.031953f
C3402 XA0.CP0 D<6> 0.238847f
C3403 XA1.CP0 D<7> 6.32554f
C3404 XA2.CP0 CK_SAMPLE 0.054172f
C3405 a_8462_2974# XB1.XA2.MP0.G 0.098184f
C3406 XA7.XA1.XA4.MP1.S AVDD 0.105303f
C3407 XA4.XA1.XA4.MP2.S EN 0.027192f
C3408 a_12422_49804# a_12422_49452# 0.010937f
C3409 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES1A.B 0.022835f
C3410 XDAC2.XC64b<1>.XRES8.B XDAC2.XC64b<1>.XRES16.B 0.1057f
C3411 XA2.CN0 XA2.XA1.XA4.LCK_N 0.012683f
C3412 XA2.XA1.CHL_OP a_4862_44348# 0.088002f
C3413 XB2.XA4.GNG m3_23150_120# 0.024512f
C3414 XB2.XA3.B m3_16526_2200# 0.024512f
C3415 XA4.CEIN VREF 0.018904f
C3416 a_21134_48572# a_21134_48220# 0.010937f
C3417 XDAC1.XC64a<0>.XRES16.B XDAC1.XC64a<0>.XRES1A.B 0.467299f
C3418 XA8.CEO CK_SAMPLE 0.025863f
C3419 XA0.CMP_OP XA2.XA1.XA4.MN2.S 0.025128f
C3420 a_3494_40828# XA1.XA1.XA1.MP3.G 0.066018f
C3421 XA0.CP1 AVDD 1.59889f
C3422 a_19982_46988# CK_SAMPLE 0.078919f
C3423 XA20.XA1.CKN a_23654_47164# 0.087851f
C3424 a_7382_47340# XA4.EN 0.071277f
C3425 XA2.XA1.XA5.MP2.S EN 0.044228f
C3426 XA5.ENO XA0.CMP_OP 0.820808f
C3427 XA8.ENO XA8.XA2.A 0.090222f
C3428 XA3.XA10.Y a_7382_48572# 0.089492f
C3429 XA8.XA10.Y XA8.XA11.MP1.S 0.010335f
C3430 XA7.ENO XA7.XA1.XA1.MP2.S 0.155821f
C3431 XA6.ENO XA7.XA1.XA1.MN2.S 0.038148f
C3432 XA1.ENO a_2342_40124# 0.024578f
C3433 XA0.CMP_OP XA0.XA1.XA4.LCK_N 0.375025f
C3434 XA0.CMP_ON XA6.XA1.XA4.LCK_N 0.276413f
C3435 XA0.XA6.Y a_n178_46988# 0.047651f
C3436 XA8.XA6.Y VREF 0.077752f
C3437 XA4.XA1.XA1.MN2.S a_9902_39772# 0.036993f
C3438 XA8.XA1.XA1.MP2.S a_21134_40124# 0.04865f
C3439 XA0.CMP_ON D<6> 0.055536f
C3440 XA1.CN1 EN 0.097358f
C3441 XA8.XA8.A a_21134_47692# 0.133834f
C3442 XA20.XA10.A a_23654_47692# 0.034262f
C3443 XA6.XA6.Y XA6.DONE 0.014904f
C3444 XA2.CN1 D<8> 0.711315f
C3445 XA3.CN1 VREF 0.618402f
C3446 XB1.XA4.GNG a_8462_1390# 0.017291f
C3447 XA1.ENO XA2.XA1.CHL_OP 0.129613f
C3448 a_11054_40476# AVDD 0.362177f
C3449 XB1.TIE_L XB1.XA1.Y 0.047823f
C3450 XA0.CEO XB1.TIE_L 0.036144f
C3451 XA4.CEO a_12422_49100# 0.07472f
C3452 XA4.XA11.Y a_11054_49100# 0.091063f
C3453 XA6.CN1 a_16094_43468# 0.070763f
C3454 XA2.ENO a_6014_40828# 0.075865f
C3455 XA8.ENO a_21134_41180# 0.072087f
C3456 XDAC2.XC64b<1>.XRES1B.B SARN 3.63755f
C3457 XA20.XA10.B CK_SAMPLE 0.176901f
C3458 a_974_48220# AVDD 0.41338f
C3459 XA0.CMP_OP XA1.XA1.XA1.MP3.G 0.142956f
C3460 XA4.XA1.XA1.MP3.S XA4.XA1.XA1.MP2.S 0.050207f
C3461 XA0.CP0 D<7> 3.31132f
C3462 XA3.CP0 AVDD 2.17073f
C3463 a_11054_46108# VREF 0.031953f
C3464 a_16094_46108# D<2> 0.011483f
C3465 XA1.CP0 CK_SAMPLE 0.054325f
C3466 XA4.ENO XA4.CN0 0.097273f
C3467 XB2.XA4.GNG m3_16598_280# 0.0666f
C3468 XA2.ENO a_8534_41884# 0.073155f
C3469 XB2.XA3.B m3_23222_3000# 0.172147f
C3470 XA8.XA11.Y AVDD 0.713612f
C3471 XA2.XA11.Y VREF 0.015286f
C3472 XA4.XA10.A a_11054_48220# 0.070424f
C3473 XA8.CEO DONE 0.093409f
C3474 XA5.XA1.XA5.MP2.S XA5.XA1.XA5.MP1.S 0.050207f
C3475 XA0.CMP_OP XA1.XA1.XA4.MN2.S 0.026188f
C3476 a_2342_40828# XA1.XA1.XA1.MP3.G 0.071498f
C3477 a_21134_46988# AVDD 0.394081f
C3478 a_12422_46988# D<3> 0.070283f
C3479 a_18614_46988# CK_SAMPLE 0.068905f
C3480 a_19982_39772# a_19982_39420# 0.010937f
C3481 XA5.XA6.Y XA5.XA6.MP3.S 0.055045f
C3482 XA2.XA1.XA4.LCK_N EN 0.038188f
C3483 XA4.XA1.XA5.MP1.S AVDD 0.102822f
C3484 XA20.XA1.CKN a_22502_47164# 0.070726f
C3485 a_7382_39420# AVDD 0.470715f
C3486 XA0.ENO a_3494_42588# 0.06916f
C3487 XA4.ENO XA0.CMP_OP 0.6934f
C3488 XA7.ENO XA8.XA2.A 0.04064f
C3489 a_12422_39772# EN 0.073293f
C3490 a_21134_46108# XA8.CP0 0.066018f
C3491 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES8.B 0.477132f
C3492 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES2.B 0.015267f
C3493 XA7.XA1.CHL_OP a_18614_41884# 0.040867f
C3494 XA1.XA1.CHL_OP XA1.XA1.XA4.MP2.S 0.050207f
C3495 XA0.CMP_ON XA5.XA1.XA5.MN1.S 0.011178f
C3496 XA0.CMP_OP a_21134_40124# 0.068085f
C3497 XA7.XA1.XA4.MN2.S XA7.XA1.XA4.MN1.S 0.050207f
C3498 a_7382_47692# AVDD 0.395235f
C3499 XA0.CMP_ON D<7> 0.056276f
C3500 XA6.CN1 D<2> 0.622769f
C3501 XA8.XA8.A a_19982_47692# 0.160931f
C3502 XA1.CN1 D<8> 0.907409f
C3503 XA2.CN1 VREF 0.618337f
C3504 a_2342_43468# AVDD 0.377891f
C3505 XA3.CN1 SARN 0.092149f
C3506 XA6.XA1.XA1.MP3.G EN 0.145483f
C3507 XA1.ENO XA1.XA1.CHL_OP 0.118011f
C3508 XA0.CP1 XA3.CP0 0.100191f
C3509 XA2.CN0 a_6014_46108# 0.103403f
C3510 XA4.CEO a_11054_49100# 0.015625f
C3511 XA4.XA11.Y a_9902_49100# 0.10248f
C3512 XDAC1.XC0.XRES1A.B SARP 3.63804f
C3513 XA6.CN1 a_14942_43468# 0.107905f
C3514 XA5.XA1.CHL_OP a_13574_42588# 0.01727f
C3515 XA2.ENO a_4862_40828# 0.132757f
C3516 XA8.ENO a_19982_41180# 0.068502f
C3517 XA20.XA10.B DONE 0.054936f
C3518 XDAC2.XC64a<0>.XRES4.B SARN 13.9307f
C3519 XA0.CMP_OP XA0.XA1.XA1.MP3.S 0.010682f
C3520 XA4.XA1.XA1.MP3.G XA4.XA1.XA1.MP2.S 0.064105f
C3521 XA2.CP0 AVDD 2.16169f
C3522 XA0.CP0 CK_SAMPLE 0.054172f
C3523 a_9614_3326# a_9614_2974# 0.010937f
C3524 XA3.XA1.XA4.MP1.S EN 0.027192f
C3525 a_11054_49804# a_11054_49452# 0.010937f
C3526 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES1A.B 0.022835f
C3527 XDAC1.XC64b<1>.XRES8.B XDAC1.XC64b<1>.XRES16.B 0.1057f
C3528 XA1.XA1.CHL_OP a_3494_44348# 0.089573f
C3529 XB2.XA4.GNG m3_16526_280# 0.105547f
C3530 XA7.XA1.CHL_OP XA8.XA1.CHL_OP 0.082663f
C3531 XB2.XA3.B m3_23150_3000# 0.0666f
C3532 a_11054_2094# SARN 0.044957f
C3533 XB1.XA1.Y SAR_IP 0.023477f
C3534 XA8.CEO AVDD 1.77861f
C3535 XA2.CEO VREF 0.367402f
C3536 a_19982_48572# a_19982_48220# 0.010937f
C3537 XA4.XA10.A a_9902_48220# 0.132671f
C3538 XDAC2.XC64a<0>.XRES2.B XDAC2.XC64a<0>.XRES1A.B 0.015267f
C3539 XA0.CMP_OP XA0.XA1.XA4.MP1.S 0.010745f
C3540 a_6014_47340# XA2.ENO 0.069707f
C3541 a_6014_39420# AVDD 0.471851f
C3542 XA4.EN XA0.CMP_OP 0.820808f
C3543 XA7.ENO XA7.XA2.A 0.090222f
C3544 a_11054_39772# EN 0.071722f
C3545 a_19982_46108# XA8.CP0 0.067789f
C3546 XA6.CN0 XA6.XA1.CHL_OP 0.037542f
C3547 XA6.ENO XA6.XA1.XA1.MP2.S 0.150467f
C3548 XA0.ENO a_974_40124# 0.025674f
C3549 XA7.XA1.CHL_OP a_17462_41884# 0.023777f
C3550 XA0.CMP_OP a_19982_40124# 0.072303f
C3551 a_6014_47692# AVDD 0.395235f
C3552 XA8.XA6.Y D<0> 0.039807f
C3553 XA7.XA8.A VREF 0.028938f
C3554 XA8.XA1.XA1.MP3.G a_21134_39420# 0.03422f
C3555 XA3.XA1.XA1.MN2.S a_8534_39772# 0.036993f
C3556 XA8.XA1.XA1.MN2.S a_19982_40124# 0.056787f
C3557 XA2.XA8.A a_6014_47340# 0.091063f
C3558 XA1.CN1 VREF 0.618402f
C3559 a_974_43468# AVDD 0.377891f
C3560 XA2.CN1 SARN 0.086984f
C3561 XB1.M1.G a_11054_1390# 0.068974f
C3562 XB2.M1.G XB2.XA4.GNG 0.250687f
C3563 XA0.ENO XA1.XA1.CHL_OP 0.13041f
C3564 XA0.CP1 XA2.CP0 0.101237f
C3565 a_21134_49452# a_21134_49100# 0.010937f
C3566 XDAC2.X16ab.XRES1A.B XDAC2.XC128b<2>.XRES1B.B 0.62895f
C3567 XA8.XA10.A DONE 0.056481f
C3568 XA20.XA10.B AVDD 1.1295f
C3569 XDAC1.XC64a<0>.XRES1B.B SARP 3.63755f
C3570 XA0.CMP_OP XA0.XA1.XA1.MP3.G 0.142977f
C3571 a_18614_48220# XA7.XA6.Y 0.071154f
C3572 XA4.XA1.XA1.MP3.G XA4.XA1.XA1.MN2.S 0.078539f
C3573 XA1.CP0 AVDD 2.17073f
C3574 XA6.XA1.XA4.MP1.S AVDD 0.105303f
C3575 XA20.XA1.CKN XA20.XA4.MP0.S 0.107674f
C3576 XB1.CKN AVDD 2.35133f
C3577 XA1.XA1.CHL_OP a_2342_44348# 0.066439f
C3578 XB2.XA4.GNG m3_23222_1080# 0.049023f
C3579 XB2.XA3.B m3_16598_3160# 0.024512f
C3580 XA7.XA11.Y AVDD 0.708074f
C3581 XA1.XA11.Y VREF 0.015777f
C3582 XA0.CMP_OP XA0.XA1.XA4.MN1.S 0.024389f
C3583 XA0.XA6.Y a_974_46108# 0.023316f
C3584 a_11054_46988# D<4> 0.068712f
C3585 a_18614_39772# a_18614_39420# 0.010937f
C3586 XA5.XA1.XA5.MP2.S AVDD 0.038567f
C3587 a_4862_47340# XA2.ENO 0.067588f
C3588 XA1.XA1.XA5.MP1.S EN 0.03516f
C3589 XA3.XA1.XA4.LCK_N D<5> 0.01587f
C3590 XA2.ENO XA0.CMP_OP 0.6934f
C3591 XA6.ENO XA7.XA2.A 0.041437f
C3592 XA2.CP0 XA3.CP0 0.959747f
C3593 XDAC2.XC128a<1>.XRES16.B XDAC2.XC32a<0>.XRES16.B 0.010386f
C3594 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES8.B 0.029725f
C3595 XA6.ENO XA6.XA1.XA1.MN2.S 0.040976f
C3596 XA2.XA2.A XA2.XA1.XA5.MN2.S 0.050207f
C3597 XA3.CN0 XA3.XA1.XA1.MP3.G 0.013311f
C3598 XA0.XA1.CHL_OP XA0.XA1.XA4.MP2.S 0.050207f
C3599 XA0.CMP_ON XA5.XA1.XA4.LCK_N 0.284482f
C3600 XA0.CMP_OP a_18614_40124# 0.073806f
C3601 XA7.XA6.Y VREF 0.078171f
C3602 XA8.XA1.XA1.MP3.G a_19982_39420# 0.023111f
C3603 XA2.XA8.A a_4862_47340# 0.127528f
C3604 a_21134_44348# VREF 0.059517f
C3605 XA5.CN1 D<3> 0.62381f
C3606 XA5.XA8.A XA5.DONE 0.1303f
C3607 XA3.CN1 D<1> 0.070704f
C3608 XA1.CN1 SARN 0.141421f
C3609 XB2.M1.G XB2.CKN 0.41624f
C3610 a_15014_1918# XB2.XA4.GNG 0.01152f
C3611 XA5.XA1.XA1.MP3.G EN 0.145483f
C3612 XA0.ENO XA0.XA1.CHL_OP 0.117946f
C3613 a_7382_40476# AVDD 0.362093f
C3614 XA5.CN0 XA7.CN0 0.364536f
C3615 XA0.CP1 XA1.CP0 0.010089f
C3616 XB1.TIE_L a_12422_2446# 0.161602f
C3617 XA4.CEIN a_11054_49100# 0.066018f
C3618 XA8.CEO XA8.XA11.Y 0.141385f
C3619 XA5.CN1 a_13574_43468# 0.109463f
C3620 XA1.ENO a_3494_40828# 0.135353f
C3621 XA7.ENO a_18614_41180# 0.06753f
C3622 XA8.XA10.A AVDD 0.769259f
C3623 a_17462_48220# XA7.XA6.Y 0.067588f
C3624 XA8.XA1.XA1.MP3.S a_21134_40476# 0.04865f
C3625 XA0.CP0 AVDD 2.16175f
C3626 a_7382_46108# VREF 0.031953f
C3627 a_19982_46108# CK_SAMPLE 0.070868f
C3628 a_8462_3326# a_8462_2974# 0.010937f
C3629 a_9902_49804# a_9902_49452# 0.010937f
C3630 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES16.B 0.063821f
C3631 XDAC2.XC64b<1>.XRES8.B XDAC2.XC64b<1>.XRES2.B 0.446669f
C3632 XB1.XA4.GNG AVDD 2.51656f
C3633 XB2.XA4.GNG m3_23150_1080# 0.024512f
C3634 XB2.XA3.B m3_16526_3160# 0.024512f
C3635 a_12422_2446# SAR_IN 0.053744f
C3636 a_18614_48572# a_18614_48220# 0.010937f
C3637 XA3.XA10.A a_8534_48220# 0.134161f
C3638 XA7.CEO AVDD 1.05093f
C3639 XA1.CEO VREF 0.018904f
C3640 XDAC1.XC64a<0>.XRES2.B XDAC1.XC64a<0>.XRES1A.B 0.015267f
C3641 XA0.CMP_OP XA1.XA1.XA4.MP2.S 0.026257f
C3642 a_974_40828# XA0.XA1.XA1.MP3.G 0.069927f
C3643 XA20.XA1.CK SARP 0.523123f
C3644 a_17462_46988# AVDD 0.395571f
C3645 a_14942_46988# CK_SAMPLE 0.070402f
C3646 XA4.XA1.XA5.MP2.S AVDD 0.038567f
C3647 XA1.XA1.XA4.LCK_N EN 0.038188f
C3648 XA1.CN0 XA3.CN1 0.418529f
C3649 XA1.ENO XA0.CMP_OP 0.820808f
C3650 XA6.ENO XA6.XA2.A 0.090222f
C3651 a_18614_46108# XA7.CP0 0.066219f
C3652 XA1.CP0 XA3.CP0 0.809357f
C3653 XA2.XA10.Y a_6014_48572# 0.091063f
C3654 XA7.XA11.MP1.S XA7.XA10.Y 0.010335f
C3655 XA5.ENO XA6.XA1.XA1.MN2.S 0.030034f
C3656 XDAC1.XC128b<2>.XRES16.B SARP 55.2956f
C3657 XA6.XA1.CHL_OP a_16094_41884# 0.023777f
C3658 XA0.XA1.CHL_OP XA0.XA1.XA4.MN2.S 0.062799f
C3659 XA0.CMP_OP a_17462_40124# 0.066394f
C3660 XA6.XA8.A VREF 0.028938f
C3661 XA7.XA1.XA1.MN2.S a_18614_40124# 0.056787f
C3662 XA2.CN1 D<1> 0.070327f
C3663 XA3.CN1 D<2> 0.065873f
C3664 XA0.CMP_ON AVDD 8.24092f
C3665 XA5.XA6.Y XA5.DONE 0.014904f
C3666 XA8.XA6.Y a_19982_47692# 0.017683f
C3667 XB2.M1.G XB2.XA4.MN1.S 0.101001f
C3668 XB1.M1.G a_8462_1390# 0.034677f
C3669 XA0.CP1 XA0.CP0 9.093941f
C3670 a_6014_40476# AVDD 0.362177f
C3671 XA7.XA1.XA1.MP3.G D<1> 0.018094f
C3672 XB1.TIE_L a_11054_2446# 0.161191f
C3673 a_19982_49452# a_19982_49100# 0.010937f
C3674 XA4.CEIN a_9902_49100# 0.070731f
C3675 XA3.XA11.Y a_8534_49100# 0.104051f
C3676 XDAC1.X16ab.XRES1A.B XDAC1.XC128b<2>.XRES1B.B 0.62895f
C3677 XDAC2.XC0.XRES1A.B SARN 3.63804f
C3678 XA5.CN1 a_12422_43468# 0.069193f
C3679 XA1.ENO a_2342_40828# 0.073834f
C3680 XA7.ENO a_17462_41180# 0.073535f
C3681 XA7.XA10.A AVDD 0.769259f
C3682 XA6.XA1.XA4.LCK_N XA6.XA1.XA4.MN2.S 0.030434f
C3683 XA8.XA1.XA1.MP3.G a_21134_40476# 0.098305f
C3684 a_21134_46108# AVDD 0.379752f
C3685 a_6014_46108# VREF 0.031953f
C3686 a_12422_46108# D<3> 0.011483f
C3687 a_18614_46108# CK_SAMPLE 0.07476f
C3688 XA7.XA1.XA4.MP2.S AVDD 0.035519f
C3689 XA2.XA1.XA4.MP1.S EN 0.027192f
C3690 XB2.M1.G AVDD 0.666052f
C3691 XA0.XA1.CHL_OP a_974_44348# 0.06801f
C3692 XB2.XA4.GNG m3_16598_1240# 0.0666f
C3693 XA1.ENO a_4862_41884# 0.074595f
C3694 XB2.XA3.B m3_23222_3960# 0.172147f
C3695 XA3.XA10.A a_7382_48220# 0.068853f
C3696 XA6.XA11.Y AVDD 0.712901f
C3697 XA0.XA11.Y VREF 0.015286f
C3698 XA0.XA1.XA4.LCK_N a_n178_41884# 0.031412f
C3699 XA0.CMP_OP XA0.XA1.XA4.MP2.S 0.026117f
C3700 a_n178_40828# XA0.XA1.XA1.MP3.G 0.067588f
C3701 a_13574_46988# CK_SAMPLE 0.068905f
C3702 XA1.CP0 XDAC1.XC64a<0>.XRES16.B 0.025998f
C3703 a_16094_46988# AVDD 0.395571f
C3704 a_17462_39772# a_17462_39420# 0.010937f
C3705 a_3494_47340# XA1.ENO 0.066018f
C3706 XA2.XA1.XA5.MN2.S EN 0.016689f
C3707 XA4.XA6.Y XA4.XA6.MP3.S 0.055045f
C3708 XA3.XA6.Y XA3.XA6.MN1.S 0.026506f
C3709 XA4.XA1.XA4.LCK_N AVDD 0.271451f
C3710 XA1.CN0 XA2.CN1 5.88308f
C3711 a_2342_39420# AVDD 0.470715f
C3712 XA0.CP1 XA0.CMP_ON 0.055536f
C3713 XA0.ENO XA0.CMP_OP 0.6934f
C3714 XA5.ENO XA6.XA2.A 0.04064f
C3715 a_7382_39772# EN 0.073293f
C3716 a_17462_46108# XA7.CP0 0.067588f
C3717 XA0.CP0 XA3.CP0 0.21972f
C3718 XA1.CP0 XA2.CP0 0.631104f
C3719 XA2.XA10.Y a_4862_48572# 0.13253f
C3720 XA8.CEO XA20.XA10.B 0.13163f
C3721 XDAC1.XC128a<1>.XRES16.B XDAC1.XC32a<0>.XRES16.B 0.010386f
C3722 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES8.B 0.029725f
C3723 XA5.ENO XA5.XA1.XA1.MN2.S 0.104122f
C3724 XA1.XA2.A XA1.XA1.XA5.MN2.S 0.050207f
C3725 XA8.XA2.A a_21134_42588# 0.129098f
C3726 XA6.XA1.CHL_OP a_14942_41884# 0.040867f
C3727 XA0.CMP_OP a_16094_40124# 0.067964f
C3728 XA7.XA1.XA4.MP2.S XA7.XA1.XA4.MP1.S 0.050207f
C3729 a_2342_47692# AVDD 0.395235f
C3730 XA2.XA6.Y a_4862_47340# 0.011912f
C3731 XA1.CN1 D<1> 0.076935f
C3732 XA2.CN1 D<2> 0.065888f
C3733 XA3.CN1 D<3> 0.065888f
C3734 a_21134_44348# D<0> 0.02026f
C3735 XA4.CN1 D<4> 0.622769f
C3736 XB1.CKN XB1.XA4.MN1.S 0.011708f
C3737 XA4.XA1.XA1.MP3.G EN 0.145483f
C3738 XA7.CEO XA8.XA11.Y 0.220689f
C3739 XA3.XA11.Y a_7382_49100# 0.089492f
C3740 XDAC1.XC0.XRES16.B SARP 55.2956f
C3741 XA4.XA1.CHL_OP a_9902_42588# 0.01727f
C3742 XA6.XA10.A AVDD 0.769259f
C3743 XDAC2.XC64a<0>.XRES1B.B SARN 3.63755f
C3744 XA2.XA1.XA4.LCK_N a_6014_41180# 0.023475f
C3745 XA5.XA1.XA4.LCK_N XA5.XA1.XA4.MN1.S 0.030434f
C3746 XA8.XA1.XA1.MP3.G a_19982_40476# 0.066018f
C3747 XA3.XA1.XA1.MP3.G XA3.XA1.XA1.MN2.S 0.078539f
C3748 XA3.XA1.XA1.MP3.S XA3.XA1.XA1.MP2.S 0.050207f
C3749 XA6.XA1.XA4.MP2.S AVDD 0.035519f
C3750 a_8534_49804# a_8534_49452# 0.010937f
C3751 XDAC1.XC64b<1>.XRES8.B XDAC1.XC64b<1>.XRES2.B 0.446669f
C3752 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES16.B 0.063821f
C3753 a_15014_1918# AVDD 0.413849f
C3754 XA0.XA1.CHL_OP a_n178_44348# 0.088002f
C3755 XB2.XA4.GNG m3_16526_1240# 0.105547f
C3756 XA5.XA1.CHL_OP XA6.XA1.CHL_OP 0.082663f
C3757 XB2.XA3.B m3_23150_3960# 0.0666f
C3758 XA3.CP0 XA0.CMP_ON 0.056088f
C3759 a_11054_2446# SAR_IP 0.053744f
C3760 a_12422_2446# SARP 0.048106f
C3761 a_17462_48572# a_17462_48220# 0.010937f
C3762 XA6.CEO AVDD 1.98375f
C3763 XA0.CEO VREF 0.367402f
C3764 XDAC2.XC64a<0>.XRES8.B XDAC2.XC64a<0>.XRES1A.B 0.029729f
C3765 XDAC2.XC64a<0>.XRES2.B XDAC2.XC64a<0>.XRES16.B 0.470901f
C3766 XA4.XA1.XA5.MP2.S XA4.XA1.XA5.MP1.S 0.050207f
C3767 XA0.CMP_OP XA0.XA1.XA4.MN2.S 0.025128f
C3768 a_2342_47340# XA1.ENO 0.071277f
C3769 XA3.XA6.Y XA3.XA6.MP1.S 0.055045f
C3770 XA1.XA1.XA5.MN2.S EN 0.016683f
C3771 XA1.CN0 XA1.CN1 2.51429f
C3772 a_974_39420# AVDD 0.471851f
C3773 XA5.ENO XA5.XA2.A 0.090222f
C3774 a_6014_39772# EN 0.071722f
C3775 XA0.CP0 XA2.CP0 0.219571f
C3776 XA5.ENO XA5.XA1.XA1.MP2.S 0.155821f
C3777 XA4.ENO XA5.XA1.XA1.MN2.S 0.038148f
C3778 XA8.XA2.A a_19982_42588# 0.089492f
C3779 XA20.XA2.VMR XA20.XA2.N2 0.025253f
C3780 XA0.CMP_OP a_14942_40124# 0.072221f
C3781 XA7.XA6.Y D<1> 0.039903f
C3782 XA6.XA6.Y VREF 0.078171f
C3783 XA20.XA11.MP1.S CK_SAMPLE 0.01103f
C3784 a_974_47692# AVDD 0.395235f
C3785 XA7.XA1.XA1.MP3.G a_18614_39420# 0.023111f
C3786 XA7.XA1.XA1.MP2.S a_17462_40124# 0.04865f
C3787 XA4.XA8.A XA4.DONE 0.1303f
C3788 a_22502_43996# AVDD 0.413321f
C3789 a_17462_44348# VREF 0.059568f
C3790 XA1.CN1 D<2> 0.104749f
C3791 XA2.CN1 D<3> 0.066027f
C3792 XA3.CN1 D<4> 0.249488f
C3793 XA5.CN0 XA6.CN0 6.33784f
C3794 XB1.TIE_L a_13862_2622# 0.011647f
C3795 XA4.CN0 XA7.CN0 0.186654f
C3796 a_18614_49452# a_18614_49100# 0.010937f
C3797 XA4.CN1 a_11054_43468# 0.070763f
C3798 XDAC2.XC0.XRES16.B D<8> 0.031495f
C3799 XA6.ENO a_16094_41180# 0.072087f
C3800 XA0.ENO a_974_40828# 0.075865f
C3801 XA5.XA10.A AVDD 0.769259f
C3802 XDAC1.XC32a<0>.XRES1A.B SARP 3.63804f
C3803 XA0.CMP_OP a_19982_40828# 0.014959f
C3804 XA2.XA1.XA4.LCK_N a_4862_41180# 0.060353f
C3805 XA3.XA1.XA1.MP3.G XA3.XA1.XA1.MP2.S 0.064105f
C3806 a_11054_46108# D<4> 0.011483f
C3807 XA3.XA1.XA4.MP2.S EN 0.027192f
C3808 XB2.XA3.B m3_16598_4120# 0.024512f
C3809 XB2.XA4.GNG m3_23222_2040# 0.049023f
C3810 XA0.ENO a_3494_41884# 0.073155f
C3811 XA7.CN0 XA0.CMP_OP 0.063388f
C3812 XA2.CP0 XA0.CMP_ON 0.057245f
C3813 XA2.XA10.A a_6014_48220# 0.070424f
C3814 XA5.XA11.Y AVDD 0.708074f
C3815 XA20.XA1.CK VREF 0.02151f
C3816 a_7382_46988# D<5> 0.070283f
C3817 a_16094_39772# a_16094_39420# 0.010937f
C3818 XA0.XA1.XA5.MP1.S EN 0.03516f
C3819 XA3.XA1.XA5.MP1.S AVDD 0.102822f
C3820 XA4.ENO XA5.XA2.A 0.041437f
C3821 XA0.CP0 XA1.CP0 4.95567f
C3822 a_16094_46108# XA6.CP0 0.066018f
C3823 XA0.CN0 XA3.CN1 0.530218f
C3824 XA1.XA10.Y a_3494_48572# 0.13402f
C3825 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES4.B 0.430615f
C3826 XDAC2.XC128b<2>.XRES16.B SARN 55.2956f
C3827 XA5.XA1.CHL_OP a_13574_41884# 0.040867f
C3828 XA20.XA2.CO XA20.XA2.N2 0.126354f
C3829 XA0.CMP_ON XA4.XA1.XA5.MN1.S 0.011062f
C3830 XA0.CMP_OP a_13574_40124# 0.073806f
C3831 XA20.XA11.MP1.S DONE 0.011819f
C3832 XA8.XA8.A CK_SAMPLE 0.02837f
C3833 XA7.XA1.XA1.MP3.G a_17462_39420# 0.03422f
C3834 a_974_49804# a_974_49452# 0.010937f
C3835 XA7.XA8.A a_18614_47692# 0.160931f
C3836 XA8.CN1 AVDD 2.03336f
C3837 a_16094_44348# VREF 0.059568f
C3838 XA1.CN1 D<3> 0.221986f
C3839 XA2.CN1 D<4> 0.06615f
C3840 XA3.CN1 D<5> 1.26542f
C3841 XB1.XA4.GNG XB1.CKN 0.142777f
C3842 XA3.XA1.XA1.MP3.G EN 0.145483f
C3843 XB1.TIE_L a_9614_2622# 0.011647f
C3844 XA6.XA1.XA1.MP3.G D<2> 0.021669f
C3845 a_2342_40476# AVDD 0.362093f
C3846 XA2.CEO a_8534_49100# 0.0733f
C3847 XA7.CEO XA7.XA11.Y 0.377598f
C3848 XA4.CN1 a_9902_43468# 0.107905f
C3849 XA3.XA1.CHL_OP a_8534_42588# 0.01727f
C3850 XA6.ENO a_14942_41180# 0.068502f
C3851 XA0.ENO a_n178_40828# 0.132757f
C3852 XA4.XA10.A AVDD 0.769259f
C3853 XA0.CMP_OP a_18614_40828# 0.014652f
C3854 a_16094_48220# XA6.XA6.Y 0.066018f
C3855 a_17462_46108# AVDD 0.378183f
C3856 a_2342_46108# VREF 0.031953f
C3857 a_14942_46108# CK_SAMPLE 0.073189f
C3858 XA5.XA1.XA4.MP1.S AVDD 0.105303f
C3859 XA2.XA1.XA4.MP2.S EN 0.027192f
C3860 a_7382_49804# a_7382_49452# 0.010937f
C3861 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES16.B 0.05157f
C3862 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES2.B 0.033713f
C3863 XB2.XA3.B m3_16526_4120# 0.024512f
C3864 XB2.XA4.GNG m3_23150_2040# 0.024512f
C3865 XA8.ENO XA8.XA1.XA4.LCK_N 0.152052f
C3866 XB1.M1.G AVDD 0.666052f
C3867 XA1.CP0 XA0.CMP_ON 0.056088f
C3868 XA20.XA2.VMR XA20.XA2.N1 0.290432f
C3869 a_16094_48572# a_16094_48220# 0.010937f
C3870 XA2.XA10.A a_4862_48220# 0.132671f
C3871 XA5.CEO AVDD 1.04893f
C3872 XDAC1.XC64a<0>.XRES8.B XDAC1.XC64a<0>.XRES1A.B 0.029729f
C3873 XDAC1.XC64a<0>.XRES2.B XDAC1.XC64a<0>.XRES16.B 0.470901f
C3874 XA4.XA1.XA4.LCK_N XA4.XA1.XA5.MN1.S 0.030434f
C3875 a_9902_46988# CK_SAMPLE 0.070402f
C3876 XA20.XA1.CK SARN 0.644014f
C3877 a_12422_46988# AVDD 0.395571f
C3878 XA8.ENO EN 0.729752f
C3879 a_974_47340# XA0.ENO 0.069707f
C3880 XA3.XA1.XA4.LCK_N AVDD 0.271288f
C3881 XA4.ENO XA4.XA2.A 0.090222f
C3882 a_14942_46108# XA6.CP0 0.067789f
C3883 XA0.CN0 XA2.CN1 0.172458f
C3884 a_21134_39772# AVDD 0.383541f
C3885 XA1.XA10.Y a_2342_48572# 0.089492f
C3886 XA6.XA10.Y XA6.XA11.MP1.S 0.010335f
C3887 XA4.ENO XA4.XA1.XA1.MP2.S 0.150467f
C3888 XA2.CN0 XA2.XA1.XA1.MP3.G 0.017163f
C3889 XA1.XA2.A XA1.XA1.XA5.MP2.S 0.050207f
C3890 XA7.XA2.A a_18614_42588# 0.091063f
C3891 XDAC1.XC128b<2>.XRES2.B SARP 7.01089f
C3892 XA5.XA1.CHL_OP a_12422_41884# 0.023777f
C3893 XA0.CMP_OP a_12422_40124# 0.066394f
C3894 XA20.XA11.MP1.S AVDD 0.107553f
C3895 XA5.XA8.A VREF 0.028938f
C3896 XA8.XA8.A DONE 0.230043f
C3897 XA2.XA1.XA1.MN2.S a_4862_39772# 0.036993f
C3898 XA6.XA1.XA1.MP2.S a_16094_40124# 0.04865f
C3899 XA7.XA8.A a_17462_47692# 0.133834f
C3900 XA7.XA6.Y a_18614_47692# 0.017683f
C3901 XA1.XA8.A a_3494_47340# 0.129098f
C3902 XA4.XA6.Y XA4.DONE 0.014904f
C3903 XA7.CN1 AVDD 2.00317f
C3904 XA1.CN1 D<4> 0.107054f
C3905 XA2.CN1 D<5> 0.066437f
C3906 XA3.CN1 D<6> 0.142972f
C3907 a_974_40476# AVDD 0.362177f
C3908 XA2.CEO a_7382_49100# 0.07472f
C3909 XA2.XA11.Y a_6014_49100# 0.091063f
C3910 a_17462_49452# a_17462_49100# 0.010937f
C3911 XDAC2.XC0.XRES16.B SARN 55.2963f
C3912 XA20.XA2.N1 XA0.CMP_OP 0.083314f
C3913 XDAC2.XC32a<0>.XRES1A.B SARN 3.63804f
C3914 XA3.XA10.A AVDD 0.769259f
C3915 XA5.XA1.XA4.LCK_N XA5.XA1.XA4.MN2.S 0.030434f
C3916 a_14942_48220# XA6.XA6.Y 0.072725f
C3917 XA7.XA1.XA1.MP3.G a_18614_40476# 0.067588f
C3918 XA7.XA1.XA1.MP3.S a_17462_40476# 0.04865f
C3919 XA2.XA1.XA1.MP3.S XA2.XA1.XA1.MP2.S 0.050207f
C3920 a_974_46108# VREF 0.031953f
C3921 a_16094_46108# AVDD 0.378183f
C3922 a_13574_46108# CK_SAMPLE 0.07476f
C3923 XA20.XA1.CKN a_23654_46812# 0.078234f
C3924 XA8.XA6.Y XA8.CP0 0.010942f
C3925 XA4.EN XA3.CN0 0.158125f
C3926 XA0.CP0 XA0.CMP_ON 0.057245f
C3927 XA7.ENO XA8.XA1.XA4.LCK_N 0.339883f
C3928 XA20.XA2.CO XA20.XA2.N1 0.310451f
C3929 XA20.XA2.VMR XA20.XA3.N2 0.146492f
C3930 XB2.XA4.GNG m3_16598_2200# 0.0666f
C3931 XA4.XA11.Y AVDD 0.712901f
C3932 a_21134_41180# a_21134_40828# 0.010937f
C3933 a_8534_46988# CK_SAMPLE 0.068905f
C3934 a_6014_46988# D<6> 0.068712f
C3935 a_11054_46988# AVDD 0.395571f
C3936 XA7.ENO EN 0.952879f
C3937 a_14942_39772# a_14942_39420# 0.010937f
C3938 a_n178_47340# XA0.ENO 0.067588f
C3939 XA3.XA6.Y XA3.CN0 0.093605f
C3940 XA1.XA1.XA5.MP2.S EN 0.044153f
C3941 XA4.EN XA4.XA2.A 0.04064f
C3942 XA0.CN0 XA1.CN1 2.86906f
C3943 a_2342_39772# EN 0.073293f
C3944 XA7.CEO XA7.XA10.A 0.010854f
C3945 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES4.B 0.430615f
C3946 XA4.ENO XA4.XA1.XA1.MN2.S 0.040976f
C3947 XA7.XA2.A a_17462_42588# 0.127528f
C3948 XA0.CMP_OP a_11054_40124# 0.067964f
C3949 XA6.XA1.XA4.MP2.S XA6.XA1.XA4.MP1.S 0.050207f
C3950 XA8.XA8.A AVDD 1.19344f
C3951 XA5.XA6.Y VREF 0.078171f
C3952 XA20.XA10.A CK_SAMPLE 0.101861f
C3953 a_n178_49804# a_n178_49452# 0.010937f
C3954 XA1.XA8.A a_2342_47340# 0.089492f
C3955 XA1.XA6.Y a_3494_47340# 0.011912f
C3956 XA6.CN1 AVDD 2.00375f
C3957 a_17462_44348# D<1> 0.02026f
C3958 XA1.CN1 D<5> 0.228006f
C3959 XA3.CN1 D<7> 0.139055f
C3960 XA2.CN1 D<6> 1.0094f
C3961 XB2.XA1.Y XB2.CKN 0.200119f
C3962 XA4.CN0 XA6.CN0 0.364802f
C3963 XA2.XA1.XA1.MP3.G EN 0.145483f
C3964 XB1.TIE_L XB2.XA2.MP0.G 0.079806f
C3965 XA2.CEO a_6014_49100# 0.015625f
C3966 XA6.CEO XA7.XA11.Y 0.293159f
C3967 XA2.XA11.Y a_4862_49100# 0.10248f
C3968 XA3.CP0 XA3.XA1.XA4.LCK_N 0.013291f
C3969 XA3.CN1 a_8534_43468# 0.112954f
C3970 XA20.XA2.N1 a_23654_43116# 0.030757f
C3971 XA5.ENO a_13574_41180# 0.06753f
C3972 XDAC1.XC0.XRES2.B SARP 7.01089f
C3973 XA2.XA10.A AVDD 0.769259f
C3974 XA7.XA1.XA1.MP3.G a_17462_40476# 0.096735f
C3975 XA2.XA1.XA1.MP3.G XA2.XA1.XA1.MP2.S 0.064105f
C3976 XA20.XA1.CKN a_22502_46812# 0.066251f
C3977 XA2.ENO XA3.CN0 0.058697f
C3978 XA1.XA1.XA4.MP1.S EN 0.027192f
C3979 a_6014_49804# a_6014_49452# 0.010937f
C3980 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES2.B 0.033713f
C3981 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES16.B 0.05157f
C3982 XA6.CN0 XA0.CMP_OP 0.06443f
C3983 XA1.CN0 XA1.XA1.XA4.LCK_N 0.012456f
C3984 XA3.XA1.CHL_OP XA4.XA1.CHL_OP 0.082663f
C3985 XA20.XA2.CO XA20.XA3.N2 0.058669f
C3986 a_8462_1918# AVDD 0.413849f
C3987 XB2.XA4.GNG m3_16526_2200# 0.105547f
C3988 XA4.CEO AVDD 1.98375f
C3989 a_14942_48572# a_14942_48220# 0.010937f
C3990 XA1.XA10.A a_3494_48220# 0.134161f
C3991 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES1A.B 0.022835f
C3992 XDAC2.XC64a<0>.XRES8.B XDAC2.XC64a<0>.XRES16.B 0.1057f
C3993 XA8.ENO VREF 0.86729f
C3994 XA6.ENO EN 1.02916f
C3995 XA4.XA6.Y XA4.XA6.MN3.S 0.089305f
C3996 XA0.XA1.XA5.MP2.S EN 0.044297f
C3997 a_13574_46108# XA5.CP0 0.066219f
C3998 XA4.EN XA3.XA2.A 0.090222f
C3999 XA5.CN0 XA5.XA1.CHL_OP 0.037394f
C4000 a_974_39772# EN 0.071936f
C4001 XA4.EN XA4.XA1.XA1.MN2.S 0.030034f
C4002 XA0.CMP_ON XA4.XA1.XA4.LCK_N 0.276413f
C4003 XA0.XA2.A XA0.XA1.XA5.MP2.S 0.050207f
C4004 XA4.XA1.CHL_OP a_11054_41884# 0.023777f
C4005 XA0.CMP_OP a_9902_40124# 0.072221f
C4006 XA6.XA6.Y D<2> 0.039903f
C4007 XA4.XA8.A VREF 0.028938f
C4008 XA20.XA10.A DONE 0.107793f
C4009 XA8.XA6.Y CK_SAMPLE 0.281644f
C4010 XA6.XA1.XA1.MP3.G a_16094_39420# 0.03422f
C4011 XA1.XA1.XA1.MN2.S a_3494_39772# 0.036993f
C4012 XA6.XA1.XA1.MN2.S a_14942_40124# 0.056787f
C4013 XA5.CN1 AVDD 2.00317f
C4014 a_12422_44348# VREF 0.059568f
C4015 XA2.CN1 D<7> 0.14594f
C4016 XA1.CN1 D<6> 0.071041f
C4017 XB2.XA1.Y XB2.XA4.MN1.S 0.011382f
C4018 XB1.M1.G XB1.XA4.MN1.S 0.101001f
C4019 XA5.CN0 XA5.XA6.MP1.S 0.028026f
C4020 XB1.TIE_L a_12422_2798# 0.104214f
C4021 XA5.XA1.XA1.MP3.G D<3> 0.017966f
C4022 XA8.XA1.XA1.MP3.S AVDD 0.139632f
C4023 a_16094_49452# a_16094_49100# 0.010937f
C4024 XA6.CEO XA7.CEO 0.432008f
C4025 XDAC2.X16ab.XRES16.B XDAC2.X16ab.XRES1A.B 0.467299f
C4026 XA3.CN1 a_7382_43468# 0.069193f
C4027 XA8.XA1.CHL_OP XA0.CMP_OP 0.036437f
C4028 XA5.ENO a_12422_41180# 0.073535f
C4029 XA1.XA10.A AVDD 0.769259f
C4030 XDAC1.XC32a<0>.XRES16.B SARP 55.2956f
C4031 XA0.CMP_OP a_14942_40828# 0.014592f
C4032 XA1.XA1.XA4.LCK_N a_3494_41180# 0.060353f
C4033 XA1.CN1 XDAC2.XC64b<1>.XRES16.B 0.027052f
C4034 XA2.XA1.XA1.MP3.G XA2.XA1.XA1.MN2.S 0.078539f
C4035 a_7382_46108# D<5> 0.011483f
C4036 XA4.XA1.XA4.MP1.S AVDD 0.105303f
C4037 XA7.CN0 XA7.XA2.A 0.035115f
C4038 a_11054_2446# SARN 0.049641f
C4039 XB2.XA1.Y AVDD 0.45332f
C4040 XB2.XA4.GNG m3_23222_3000# 0.049023f
C4041 XB1.XA3.B m3_974_120# 0.0666f
C4042 a_12422_2798# SAR_IN 0.02841f
C4043 XA3.XA11.Y AVDD 0.708074f
C4044 XA1.XA10.A a_2342_48220# 0.068853f
C4045 a_19982_41180# a_19982_40828# 0.010937f
C4046 XA7.ENO VREF 0.879117f
C4047 XA5.ENO EN 0.952619f
C4048 a_13574_39772# a_13574_39420# 0.010937f
C4049 XA20.XA1.CKN XA20.XA10.MN1.S 0.097398f
C4050 XA2.XA1.XA5.MP1.S AVDD 0.102822f
C4051 XA2.XA1.XA4.LCK_N D<6> 0.015734f
C4052 XA0.XA1.XA4.LCK_N EN 0.37807f
C4053 a_15014_334# a_15014_n18# 0.010937f
C4054 a_12422_46108# XA5.CP0 0.067588f
C4055 XA2.ENO XA3.XA2.A 0.041437f
C4056 a_17462_39772# AVDD 0.382762f
C4057 a_n178_39772# EN 0.079159f
C4058 XA6.CEO XA7.XA10.A 0.019775f
C4059 XA4.EN XA3.XA1.XA1.MN2.S 0.104122f
C4060 XA20.XA1.CK XA20.XA1.MP0.S 0.010345f
C4061 XA0.CMP_ON XA3.XA1.XA5.MN1.S 0.011178f
C4062 XA4.XA1.CHL_OP a_9902_41884# 0.040867f
C4063 XA6.XA2.A a_16094_42588# 0.129098f
C4064 XDAC2.XC128b<2>.XRES2.B SARN 7.01089f
C4065 XA0.CMP_OP a_8534_40124# 0.073806f
C4066 XA20.XA10.A AVDD 0.660701f
C4067 XA8.XA6.Y DONE 0.03889f
C4068 XA6.XA1.XA1.MP3.G a_14942_39420# 0.023111f
C4069 XA6.XA8.A a_16094_47692# 0.133834f
C4070 XA3.XA8.A XA3.DONE 0.1303f
C4071 XA4.CN1 AVDD 2.00375f
C4072 a_11054_44348# VREF 0.059568f
C4073 a_16094_44348# D<2> 0.02026f
C4074 XA1.CN1 D<7> 1.13793f
C4075 a_15014_1918# XB2.M1.G 0.071041f
C4076 XB2.XA1.MP0.G XB2.XA4.GNG 0.018609f
C4077 XB1.M1.G XB1.CKN 0.41624f
C4078 XA1.CN0 a_2342_46108# 0.101833f
C4079 XB1.TIE_L a_11054_2798# 0.102644f
C4080 XA1.XA1.XA1.MP3.G EN 0.145483f
C4081 XA8.XA1.XA1.MP3.G AVDD 1.08373f
C4082 XA1.CEO a_6014_49100# 0.066018f
C4083 XA6.CEO XA6.XA11.Y 0.158152f
C4084 CK_SAMPLE_BSSW AVSS 23.03f
C4085 SAR_IN AVSS 1.66024f
C4086 SAR_IP AVSS 1.66009f
C4087 SARP AVSS 0.134912p
C4088 EN AVSS 7.81241f
C4089 D<8> AVSS 19.0987f
C4090 VREF AVSS 21.5694f
C4091 SARN AVSS 0.134165p
C4092 D<0> AVSS 0.887067f
C4093 D<1> AVSS 11.4543f
C4094 D<2> AVSS 8.907419f
C4095 D<3> AVSS 7.66246f
C4096 D<4> AVSS 8.376559f
C4097 D<5> AVSS 7.67676f
C4098 D<6> AVSS 8.76668f
C4099 D<7> AVSS 7.67274f
C4100 CK_SAMPLE AVSS 21.392f
C4101 DONE AVSS 1.0388f
C4102 AVDD AVSS 0.517053p
C4103 li_14960_5188# AVSS 0.039452f $ **FLOATING
C4104 li_9168_5188# AVSS 0.039452f $ **FLOATING
C4105 XDAC2.XC1.XRES1A.B AVSS 7.69832f
C4106 XDAC1.XC1.XRES1A.B AVSS 7.69832f
C4107 li_14960_5800# AVSS 0.035609f $ **FLOATING
C4108 li_9168_5800# AVSS 0.035609f $ **FLOATING
C4109 XDAC2.XC1.XRES16.B AVSS 15.4598f
C4110 XDAC1.XC1.XRES16.B AVSS 15.4598f
C4111 li_14960_6412# AVSS 0.035609f $ **FLOATING
C4112 li_9168_6412# AVSS 0.035609f $ **FLOATING
C4113 XDAC2.XC1.XRES2.B AVSS 8.084061f
C4114 XDAC1.XC1.XRES2.B AVSS 8.084061f
C4115 li_14960_7024# AVSS 0.035609f $ **FLOATING
C4116 li_9168_7024# AVSS 0.035609f $ **FLOATING
C4117 XDAC2.XC1.XRES8.B AVSS 11.2692f
C4118 XDAC1.XC1.XRES8.B AVSS 11.2692f
C4119 li_14960_7636# AVSS 0.035609f $ **FLOATING
C4120 li_9168_7636# AVSS 0.035609f $ **FLOATING
C4121 XDAC2.XC1.XRES4.B AVSS 9.198461f
C4122 XDAC1.XC1.XRES4.B AVSS 9.198461f
C4123 li_14960_8248# AVSS 0.033725f $ **FLOATING
C4124 li_9168_8248# AVSS 0.033725f $ **FLOATING
C4125 XDAC2.XC1.XRES1B.B AVSS 7.46832f
C4126 XDAC1.XC1.XRES1B.B AVSS 7.46832f
C4127 li_14960_8660# AVSS 0.033725f $ **FLOATING
C4128 li_9168_8660# AVSS 0.033725f $ **FLOATING
C4129 XDAC2.XC64a<0>.XRES1A.B AVSS 7.45743f
C4130 XDAC1.XC64a<0>.XRES1A.B AVSS 7.45743f
C4131 li_14960_9272# AVSS 0.035609f $ **FLOATING
C4132 li_9168_9272# AVSS 0.035609f $ **FLOATING
C4133 XDAC2.XC64a<0>.XRES16.B AVSS 15.4738f
C4134 XDAC1.XC64a<0>.XRES16.B AVSS 15.4738f
C4135 li_14960_9884# AVSS 0.035609f $ **FLOATING
C4136 li_9168_9884# AVSS 0.035609f $ **FLOATING
C4137 XDAC2.XC64a<0>.XRES2.B AVSS 8.08342f
C4138 XDAC1.XC64a<0>.XRES2.B AVSS 8.08342f
C4139 li_14960_10496# AVSS 0.035621f $ **FLOATING
C4140 li_9168_10496# AVSS 0.035621f $ **FLOATING
C4141 XDAC2.XC64a<0>.XRES8.B AVSS 11.2692f
C4142 XDAC1.XC64a<0>.XRES8.B AVSS 11.2692f
C4143 li_14960_11108# AVSS 0.035677f $ **FLOATING
C4144 li_9168_11108# AVSS 0.035677f $ **FLOATING
C4145 XDAC2.XC64a<0>.XRES4.B AVSS 9.198461f
C4146 XDAC1.XC64a<0>.XRES4.B AVSS 9.198461f
C4147 li_14960_11720# AVSS 0.034178f $ **FLOATING
C4148 li_9168_11720# AVSS 0.034178f $ **FLOATING
C4149 XDAC2.XC64a<0>.XRES1B.B AVSS 7.46832f
C4150 XDAC1.XC64a<0>.XRES1B.B AVSS 7.46832f
C4151 li_14960_12132# AVSS 0.037637f $ **FLOATING
C4152 XDAC2.XC32a<0>.XRES1A.B AVSS 7.45868f
C4153 li_9168_12132# AVSS 0.037637f $ **FLOATING
C4154 XDAC1.XC32a<0>.XRES1A.B AVSS 7.45868f
C4155 li_14960_12744# AVSS 0.035807f $ **FLOATING
C4156 li_9168_12744# AVSS 0.035807f $ **FLOATING
C4157 XDAC2.XC32a<0>.XRES16.B AVSS 15.474201f
C4158 XDAC1.XC32a<0>.XRES16.B AVSS 15.474201f
C4159 li_14960_13356# AVSS 0.035656f $ **FLOATING
C4160 li_9168_13356# AVSS 0.035656f $ **FLOATING
C4161 XDAC2.XC32a<0>.XRES2.B AVSS 8.08342f
C4162 XDAC1.XC32a<0>.XRES2.B AVSS 8.08342f
C4163 li_14960_13968# AVSS 0.035609f $ **FLOATING
C4164 li_9168_13968# AVSS 0.035609f $ **FLOATING
C4165 XDAC2.XC32a<0>.XRES8.B AVSS 11.2692f
C4166 XDAC1.XC32a<0>.XRES8.B AVSS 11.2692f
C4167 li_14960_14580# AVSS 0.035609f $ **FLOATING
C4168 li_9168_14580# AVSS 0.035609f $ **FLOATING
C4169 XDAC2.XC32a<0>.XRES4.B AVSS 9.198461f
C4170 XDAC1.XC32a<0>.XRES4.B AVSS 9.198461f
C4171 li_14960_15192# AVSS 0.033725f $ **FLOATING
C4172 li_9168_15192# AVSS 0.033725f $ **FLOATING
C4173 XDAC2.XC32a<0>.XRES1B.B AVSS 7.46832f
C4174 XDAC1.XC32a<0>.XRES1B.B AVSS 7.46832f
C4175 li_14960_15604# AVSS 0.033725f $ **FLOATING
C4176 li_9168_15604# AVSS 0.033725f $ **FLOATING
C4177 XDAC2.XC128a<1>.XRES1A.B AVSS 7.45743f
C4178 XDAC1.XC128a<1>.XRES1A.B AVSS 7.45743f
C4179 li_14960_16216# AVSS 0.035609f $ **FLOATING
C4180 li_9168_16216# AVSS 0.035609f $ **FLOATING
C4181 XDAC2.XC128a<1>.XRES16.B AVSS 15.470799f
C4182 XDAC1.XC128a<1>.XRES16.B AVSS 15.470799f
C4183 li_14960_16828# AVSS 0.035609f $ **FLOATING
C4184 li_9168_16828# AVSS 0.035609f $ **FLOATING
C4185 XDAC2.XC128a<1>.XRES2.B AVSS 8.08342f
C4186 XDAC1.XC128a<1>.XRES2.B AVSS 8.08342f
C4187 li_14960_17440# AVSS 0.035609f $ **FLOATING
C4188 li_9168_17440# AVSS 0.035609f $ **FLOATING
C4189 XDAC2.XC128a<1>.XRES8.B AVSS 11.2692f
C4190 XDAC1.XC128a<1>.XRES8.B AVSS 11.2692f
C4191 li_14960_18052# AVSS 0.035609f $ **FLOATING
C4192 li_9168_18052# AVSS 0.035609f $ **FLOATING
C4193 XDAC2.XC128a<1>.XRES4.B AVSS 9.198461f
C4194 XDAC1.XC128a<1>.XRES4.B AVSS 9.198461f
C4195 li_14960_18664# AVSS 0.033725f $ **FLOATING
C4196 li_9168_18664# AVSS 0.033725f $ **FLOATING
C4197 XDAC2.XC128a<1>.XRES1B.B AVSS 7.46832f
C4198 XDAC1.XC128a<1>.XRES1B.B AVSS 7.46832f
C4199 li_14960_19076# AVSS 0.033725f $ **FLOATING
C4200 li_9168_19076# AVSS 0.033725f $ **FLOATING
C4201 XDAC2.XC128b<2>.XRES1A.B AVSS 7.45743f
C4202 XDAC1.XC128b<2>.XRES1A.B AVSS 7.45743f
C4203 li_14960_19688# AVSS 0.035609f $ **FLOATING
C4204 li_9168_19688# AVSS 0.035609f $ **FLOATING
C4205 XDAC2.XC128b<2>.XRES16.B AVSS 15.471701f
C4206 XDAC1.XC128b<2>.XRES16.B AVSS 15.471701f
C4207 li_14960_20300# AVSS 0.035609f $ **FLOATING
C4208 li_9168_20300# AVSS 0.035609f $ **FLOATING
C4209 XDAC2.XC128b<2>.XRES2.B AVSS 8.08342f
C4210 XDAC1.XC128b<2>.XRES2.B AVSS 8.08342f
C4211 li_14960_20912# AVSS 0.035609f $ **FLOATING
C4212 li_9168_20912# AVSS 0.035609f $ **FLOATING
C4213 XDAC2.XC128b<2>.XRES8.B AVSS 11.2692f
C4214 XDAC1.XC128b<2>.XRES8.B AVSS 11.2692f
C4215 li_14960_21524# AVSS 0.035609f $ **FLOATING
C4216 li_9168_21524# AVSS 0.035609f $ **FLOATING
C4217 XDAC2.XC128b<2>.XRES4.B AVSS 9.198461f
C4218 XDAC1.XC128b<2>.XRES4.B AVSS 9.198461f
C4219 li_14960_22136# AVSS 0.033725f $ **FLOATING
C4220 li_9168_22136# AVSS 0.033725f $ **FLOATING
C4221 XDAC2.XC128b<2>.XRES1B.B AVSS 7.46832f
C4222 XDAC1.XC128b<2>.XRES1B.B AVSS 7.46832f
C4223 li_14960_22548# AVSS 0.033725f $ **FLOATING
C4224 li_9168_22548# AVSS 0.033725f $ **FLOATING
C4225 XDAC2.X16ab.XRES1A.B AVSS 7.45743f
C4226 XDAC1.X16ab.XRES1A.B AVSS 7.45743f
C4227 li_14960_23160# AVSS 0.035609f $ **FLOATING
C4228 li_9168_23160# AVSS 0.035609f $ **FLOATING
C4229 XDAC2.X16ab.XRES16.B AVSS 15.473901f
C4230 XDAC1.X16ab.XRES16.B AVSS 15.473901f
C4231 li_14960_23772# AVSS 0.035609f $ **FLOATING
C4232 li_9168_23772# AVSS 0.035609f $ **FLOATING
C4233 XDAC2.X16ab.XRES2.B AVSS 8.08342f
C4234 XDAC1.X16ab.XRES2.B AVSS 8.08342f
C4235 li_14960_24384# AVSS 0.035609f $ **FLOATING
C4236 li_9168_24384# AVSS 0.035609f $ **FLOATING
C4237 XDAC2.X16ab.XRES8.B AVSS 11.2692f
C4238 XDAC1.X16ab.XRES8.B AVSS 11.2692f
C4239 li_14960_24996# AVSS 0.035609f $ **FLOATING
C4240 li_9168_24996# AVSS 0.035609f $ **FLOATING
C4241 XDAC2.X16ab.XRES4.B AVSS 9.198461f
C4242 XDAC1.X16ab.XRES4.B AVSS 9.198461f
C4243 li_14960_25608# AVSS 0.033725f $ **FLOATING
C4244 li_9168_25608# AVSS 0.033725f $ **FLOATING
C4245 XDAC2.X16ab.XRES1B.B AVSS 7.46832f
C4246 XDAC1.X16ab.XRES1B.B AVSS 7.46832f
C4247 li_14960_26020# AVSS 0.033725f $ **FLOATING
C4248 li_9168_26020# AVSS 0.033725f $ **FLOATING
C4249 XDAC2.XC64b<1>.XRES1A.B AVSS 7.45743f
C4250 XDAC1.XC64b<1>.XRES1A.B AVSS 7.45743f
C4251 li_14960_26632# AVSS 0.035609f $ **FLOATING
C4252 li_9168_26632# AVSS 0.035609f $ **FLOATING
C4253 XDAC2.XC64b<1>.XRES16.B AVSS 15.472301f
C4254 XDAC1.XC64b<1>.XRES16.B AVSS 15.472301f
C4255 li_14960_27244# AVSS 0.035609f $ **FLOATING
C4256 li_9168_27244# AVSS 0.035609f $ **FLOATING
C4257 XDAC2.XC64b<1>.XRES2.B AVSS 8.08342f
C4258 XDAC1.XC64b<1>.XRES2.B AVSS 8.08342f
C4259 li_14960_27856# AVSS 0.035609f $ **FLOATING
C4260 li_9168_27856# AVSS 0.035609f $ **FLOATING
C4261 XDAC2.XC64b<1>.XRES8.B AVSS 11.2692f
C4262 XDAC1.XC64b<1>.XRES8.B AVSS 11.2692f
C4263 li_14960_28468# AVSS 0.035609f $ **FLOATING
C4264 li_9168_28468# AVSS 0.035609f $ **FLOATING
C4265 XDAC2.XC64b<1>.XRES4.B AVSS 9.198461f
C4266 XDAC1.XC64b<1>.XRES4.B AVSS 9.198461f
C4267 li_14960_29080# AVSS 0.033725f $ **FLOATING
C4268 li_9168_29080# AVSS 0.033725f $ **FLOATING
C4269 XDAC2.XC64b<1>.XRES1B.B AVSS 7.46832f
C4270 XDAC1.XC64b<1>.XRES1B.B AVSS 7.46832f
C4271 li_14960_29492# AVSS 0.033725f $ **FLOATING
C4272 li_9168_29492# AVSS 0.033725f $ **FLOATING
C4273 XDAC2.XC0.XRES1A.B AVSS 7.45743f
C4274 XDAC1.XC0.XRES1A.B AVSS 7.45743f
C4275 li_14960_30104# AVSS 0.035609f $ **FLOATING
C4276 li_9168_30104# AVSS 0.035609f $ **FLOATING
C4277 XDAC2.XC0.XRES16.B AVSS 15.470701f
C4278 XDAC1.XC0.XRES16.B AVSS 15.470701f
C4279 li_14960_30716# AVSS 0.035609f $ **FLOATING
C4280 li_9168_30716# AVSS 0.035609f $ **FLOATING
C4281 XDAC2.XC0.XRES2.B AVSS 8.08342f
C4282 XDAC1.XC0.XRES2.B AVSS 8.08342f
C4283 li_14960_31328# AVSS 0.035609f $ **FLOATING
C4284 li_9168_31328# AVSS 0.035609f $ **FLOATING
C4285 XDAC2.XC0.XRES8.B AVSS 11.2716f
C4286 XDAC1.XC0.XRES8.B AVSS 11.2716f
C4287 li_14960_31940# AVSS 0.035609f $ **FLOATING
C4288 li_9168_31940# AVSS 0.035609f $ **FLOATING
C4289 XDAC2.XC0.XRES4.B AVSS 9.20524f
C4290 XDAC1.XC0.XRES4.B AVSS 9.20524f
C4291 li_14960_32552# AVSS 0.039464f $ **FLOATING
C4292 li_9168_32552# AVSS 0.039464f $ **FLOATING
C4293 XDAC2.XC0.XRES1B.B AVSS 8.169431f
C4294 XDAC1.XC0.XRES1B.B AVSS 8.166241f
C4295 a_15014_n18# AVSS 0.097214f $ **FLOATING
C4296 a_13862_n18# AVSS 0.544578f $ **FLOATING
C4297 a_12422_n18# AVSS 0.429487f $ **FLOATING
C4298 a_11054_n18# AVSS 0.429072f $ **FLOATING
C4299 a_9614_n18# AVSS 0.545733f $ **FLOATING
C4300 a_8462_n18# AVSS 0.097214f $ **FLOATING
C4301 a_13862_334# AVSS 0.492909f $ **FLOATING
C4302 a_12422_334# AVSS 0.352975f $ **FLOATING
C4303 a_11054_334# AVSS 0.352975f $ **FLOATING
C4304 a_9614_334# AVSS 0.491371f $ **FLOATING
C4305 a_13862_686# AVSS 0.37586f $ **FLOATING
C4306 a_12422_686# AVSS 0.352702f $ **FLOATING
C4307 a_11054_686# AVSS 0.352702f $ **FLOATING
C4308 a_9614_686# AVSS 0.375878f $ **FLOATING
C4309 a_12422_1038# AVSS 0.352487f $ **FLOATING
C4310 a_11054_1038# AVSS 0.352487f $ **FLOATING
C4311 XB2.XA3.B AVSS 41.8193f
C4312 XB2.XA3.MP0.S AVSS 0.703969f
C4313 XB1.XA3.B AVSS 41.8193f
C4314 XB1.XA3.MP0.S AVSS 0.704013f
C4315 a_13862_1390# AVSS 0.397761f $ **FLOATING
C4316 a_12422_1390# AVSS 0.354407f $ **FLOATING
C4317 a_11054_1390# AVSS 0.354407f $ **FLOATING
C4318 a_9614_1390# AVSS 0.397761f $ **FLOATING
C4319 XB2.XA4.GNG AVSS 37.6698f
C4320 XB2.CKN AVSS 2.39378f
C4321 XB2.XA4.MN1.S AVSS 0.104384f
C4322 a_12422_1742# AVSS 0.352432f $ **FLOATING
C4323 a_11054_1742# AVSS 0.352432f $ **FLOATING
C4324 XB1.XA4.MN1.S AVSS 0.104384f
C4325 XB1.CKN AVSS 2.39386f
C4326 XB1.XA4.GNG AVSS 37.6698f
C4327 XB2.M1.G AVSS 3.13376f
C4328 a_13862_1918# AVSS 0.389641f $ **FLOATING
C4329 XB1.M1.G AVSS 3.09498f
C4330 a_9614_1918# AVSS 0.389641f $ **FLOATING
C4331 XB2.XA1.Y AVSS 0.975394f
C4332 a_12422_2094# AVSS 0.352456f $ **FLOATING
C4333 a_11054_2094# AVSS 0.352456f $ **FLOATING
C4334 XB2.XA1.MP0.G AVSS 0.797677f
C4335 a_13862_2270# AVSS 0.470686f $ **FLOATING
C4336 XB1.XA1.MP0.G AVSS 0.797677f
C4337 XB1.XA1.Y AVSS 0.975394f
C4338 a_9614_2270# AVSS 0.472257f $ **FLOATING
C4339 a_12422_2446# AVSS 0.353103f $ **FLOATING
C4340 a_11054_2446# AVSS 0.353103f $ **FLOATING
C4341 a_13862_2622# AVSS 0.493494f $ **FLOATING
C4342 a_9614_2622# AVSS 0.491924f $ **FLOATING
C4343 XB2.XA2.MP0.G AVSS 0.59762f
C4344 a_12422_2798# AVSS 0.433341f $ **FLOATING
C4345 a_11054_2798# AVSS 0.433756f $ **FLOATING
C4346 a_13862_2974# AVSS 0.472546f $ **FLOATING
C4347 a_15014_3326# AVSS 0.090299f $ **FLOATING
C4348 a_13862_3326# AVSS 0.542115f $ **FLOATING
C4349 XB1.XA2.MP0.G AVSS 0.59762f
C4350 a_9614_2974# AVSS 0.474117f $ **FLOATING
C4351 a_9614_3326# AVSS 0.54096f $ **FLOATING
C4352 a_8462_3326# AVSS 0.090299f $ **FLOATING
C4353 a_23654_39068# AVSS 0.532853f $ **FLOATING
C4354 a_22502_39068# AVSS 0.088967f $ **FLOATING
C4355 a_21134_39068# AVSS 0.088967f $ **FLOATING
C4356 a_19982_39068# AVSS 0.531076f $ **FLOATING
C4357 a_18614_39068# AVSS 0.532231f $ **FLOATING
C4358 a_17462_39068# AVSS 0.088807f $ **FLOATING
C4359 a_16094_39068# AVSS 0.088807f $ **FLOATING
C4360 a_14942_39068# AVSS 0.531076f $ **FLOATING
C4361 a_13574_39068# AVSS 0.532231f $ **FLOATING
C4362 a_12422_39068# AVSS 0.088807f $ **FLOATING
C4363 a_11054_39068# AVSS 0.088807f $ **FLOATING
C4364 a_9902_39068# AVSS 0.530746f $ **FLOATING
C4365 a_8534_39068# AVSS 0.531355f $ **FLOATING
C4366 a_7382_39068# AVSS 0.088807f $ **FLOATING
C4367 a_6014_39068# AVSS 0.088807f $ **FLOATING
C4368 a_4862_39068# AVSS 0.530504f $ **FLOATING
C4369 a_3494_39068# AVSS 0.531221f $ **FLOATING
C4370 a_2342_39068# AVSS 0.088807f $ **FLOATING
C4371 a_974_39068# AVSS 0.088807f $ **FLOATING
C4372 a_n178_39068# AVSS 0.532136f $ **FLOATING
C4373 a_23654_39420# AVSS 0.501428f $ **FLOATING
C4374 a_19982_39420# AVSS 0.471864f $ **FLOATING
C4375 a_18614_39420# AVSS 0.46804f $ **FLOATING
C4376 a_14942_39420# AVSS 0.471864f $ **FLOATING
C4377 a_13574_39420# AVSS 0.46804f $ **FLOATING
C4378 a_9902_39420# AVSS 0.471204f $ **FLOATING
C4379 a_8534_39420# AVSS 0.466319f $ **FLOATING
C4380 a_4862_39420# AVSS 0.47072f $ **FLOATING
C4381 a_3494_39420# AVSS 0.466051f $ **FLOATING
C4382 a_n178_39420# AVSS 0.472352f $ **FLOATING
C4383 a_19982_39772# AVSS 0.388068f $ **FLOATING
C4384 a_18614_39772# AVSS 0.386549f $ **FLOATING
C4385 a_14942_39772# AVSS 0.388068f $ **FLOATING
C4386 a_13574_39772# AVSS 0.386549f $ **FLOATING
C4387 a_9902_39772# AVSS 0.38747f $ **FLOATING
C4388 a_8534_39772# AVSS 0.384797f $ **FLOATING
C4389 a_4862_39772# AVSS 0.387164f $ **FLOATING
C4390 a_3494_39772# AVSS 0.384529f $ **FLOATING
C4391 a_n178_39772# AVSS 0.38817f $ **FLOATING
C4392 a_19982_40124# AVSS 0.371141f $ **FLOATING
C4393 a_18614_40124# AVSS 0.369092f $ **FLOATING
C4394 a_14942_40124# AVSS 0.371141f $ **FLOATING
C4395 a_13574_40124# AVSS 0.369092f $ **FLOATING
C4396 a_9902_40124# AVSS 0.37048f $ **FLOATING
C4397 a_8534_40124# AVSS 0.36734f $ **FLOATING
C4398 a_4862_40124# AVSS 0.369997f $ **FLOATING
C4399 a_3494_40124# AVSS 0.367072f $ **FLOATING
C4400 a_n178_40124# AVSS 0.371003f $ **FLOATING
C4401 XA8.XA1.XA1.MN2.S AVSS 0.514227f
C4402 XA7.XA1.XA1.MN2.S AVSS 0.482217f
C4403 XA6.XA1.XA1.MN2.S AVSS 0.506261f
C4404 XA5.XA1.XA1.MN2.S AVSS 0.482217f
C4405 XA4.XA1.XA1.MN2.S AVSS 0.506261f
C4406 XA3.XA1.XA1.MN2.S AVSS 0.482217f
C4407 XA2.XA1.XA1.MN2.S AVSS 0.506261f
C4408 XA1.XA1.XA1.MN2.S AVSS 0.482217f
C4409 XA0.XA1.XA1.MN2.S AVSS 0.506261f
C4410 XA20.XA1.MP0.S AVSS 0.614508f
C4411 a_19982_40476# AVSS 0.40664f $ **FLOATING
C4412 a_18614_40476# AVSS 0.40664f $ **FLOATING
C4413 a_14942_40476# AVSS 0.40664f $ **FLOATING
C4414 a_13574_40476# AVSS 0.40664f $ **FLOATING
C4415 a_9902_40476# AVSS 0.406071f $ **FLOATING
C4416 a_8534_40476# AVSS 0.404979f $ **FLOATING
C4417 a_4862_40476# AVSS 0.405588f $ **FLOATING
C4418 a_3494_40476# AVSS 0.404711f $ **FLOATING
C4419 a_n178_40476# AVSS 0.406594f $ **FLOATING
C4420 XA8.XA1.XA1.MP3.G AVSS 0.759935f
C4421 XA7.XA1.XA1.MP3.G AVSS 0.736475f
C4422 XA6.XA1.XA1.MP3.G AVSS 0.750304f
C4423 XA5.XA1.XA1.MP3.G AVSS 0.736475f
C4424 XA4.XA1.XA1.MP3.G AVSS 0.749258f
C4425 XA3.XA1.XA1.MP3.G AVSS 0.732153f
C4426 XA2.XA1.XA1.MP3.G AVSS 0.747923f
C4427 XA1.XA1.XA1.MP3.G AVSS 0.731542f
C4428 XA0.XA1.XA1.MP3.G AVSS 0.750694f
C4429 a_23654_40828# AVSS 0.404746f $ **FLOATING
C4430 a_19982_40828# AVSS 0.388483f $ **FLOATING
C4431 a_18614_40828# AVSS 0.388483f $ **FLOATING
C4432 a_14942_40828# AVSS 0.388483f $ **FLOATING
C4433 a_13574_40828# AVSS 0.388483f $ **FLOATING
C4434 a_9902_40828# AVSS 0.387914f $ **FLOATING
C4435 a_8534_40828# AVSS 0.386822f $ **FLOATING
C4436 a_4862_40828# AVSS 0.387431f $ **FLOATING
C4437 a_3494_40828# AVSS 0.386554f $ **FLOATING
C4438 a_n178_40828# AVSS 0.388437f $ **FLOATING
C4439 a_19982_41180# AVSS 0.395265f $ **FLOATING
C4440 a_18614_41180# AVSS 0.3953f $ **FLOATING
C4441 a_14942_41180# AVSS 0.3953f $ **FLOATING
C4442 a_13574_41180# AVSS 0.3953f $ **FLOATING
C4443 a_9902_41180# AVSS 0.394731f $ **FLOATING
C4444 a_8534_41180# AVSS 0.393639f $ **FLOATING
C4445 a_4862_41180# AVSS 0.394248f $ **FLOATING
C4446 a_3494_41180# AVSS 0.393371f $ **FLOATING
C4447 a_n178_41180# AVSS 0.395254f $ **FLOATING
C4448 XA8.XA1.XA4.MN1.S AVSS 0.084824f
C4449 XA7.XA1.XA4.MN1.S AVSS 0.098298f
C4450 XA8.XA1.XA4.MN2.S AVSS 0.03705f
C4451 XA7.XA1.XA4.MN2.S AVSS 0.026202f
C4452 XA6.XA1.XA4.MN1.S AVSS 0.098298f
C4453 XA5.XA1.XA4.MN1.S AVSS 0.098298f
C4454 XA6.XA1.XA4.MN2.S AVSS 0.026202f
C4455 XA5.XA1.XA4.MN2.S AVSS 0.026202f
C4456 XA4.XA1.XA4.MN1.S AVSS 0.098298f
C4457 XA3.XA1.XA4.MN1.S AVSS 0.098298f
C4458 XA4.XA1.XA4.MN2.S AVSS 0.026202f
C4459 XA3.XA1.XA4.MN2.S AVSS 0.026202f
C4460 XA2.XA1.XA4.MN1.S AVSS 0.098298f
C4461 XA1.XA1.XA4.MN1.S AVSS 0.098298f
C4462 XA2.XA1.XA4.MN2.S AVSS 0.026202f
C4463 XA1.XA1.XA4.MN2.S AVSS 0.026202f
C4464 XA0.XA1.XA4.MN1.S AVSS 0.098298f
C4465 XA0.XA1.XA4.MN2.S AVSS 0.026202f
C4466 XA20.XA2.N2 AVSS 0.321933f
C4467 a_19982_41884# AVSS 0.39655f $ **FLOATING
C4468 a_18614_41884# AVSS 0.396102f $ **FLOATING
C4469 a_14942_41884# AVSS 0.39663f $ **FLOATING
C4470 a_13574_41884# AVSS 0.396102f $ **FLOATING
C4471 a_9902_41884# AVSS 0.396061f $ **FLOATING
C4472 a_8534_41884# AVSS 0.394528f $ **FLOATING
C4473 a_4862_41884# AVSS 0.395577f $ **FLOATING
C4474 a_3494_41884# AVSS 0.39426f $ **FLOATING
C4475 a_n178_41884# AVSS 0.396584f $ **FLOATING
C4476 a_23654_42236# AVSS 0.40374f $ **FLOATING
C4477 XA8.XA1.XA5.MN1.S AVSS 0.08587f
C4478 XA8.XA1.XA4.LCK_N AVSS 1.27154f
C4479 XA7.XA1.XA5.MN1.S AVSS 0.10078f
C4480 XA7.XA1.XA4.LCK_N AVSS 1.26583f
C4481 XA8.XA1.XA5.MN2.S AVSS 0.044592f
C4482 XA7.XA1.XA5.MN2.S AVSS 0.049396f
C4483 XA6.XA1.XA5.MN1.S AVSS 0.10078f
C4484 XA6.XA1.XA4.LCK_N AVSS 1.26677f
C4485 XA5.XA1.XA5.MN1.S AVSS 0.10078f
C4486 XA5.XA1.XA4.LCK_N AVSS 1.26583f
C4487 XA6.XA1.XA5.MN2.S AVSS 0.049396f
C4488 XA5.XA1.XA5.MN2.S AVSS 0.049396f
C4489 XA4.XA1.XA5.MN1.S AVSS 0.10078f
C4490 XA4.XA1.XA4.LCK_N AVSS 1.26386f
C4491 XA3.XA1.XA5.MN1.S AVSS 0.10078f
C4492 XA3.XA1.XA4.LCK_N AVSS 1.25643f
C4493 XA4.XA1.XA5.MN2.S AVSS 0.049396f
C4494 XA3.XA1.XA5.MN2.S AVSS 0.049396f
C4495 XA2.XA1.XA5.MN1.S AVSS 0.10078f
C4496 XA2.XA1.XA4.LCK_N AVSS 1.26168f
C4497 XA1.XA1.XA5.MN1.S AVSS 0.10078f
C4498 XA1.XA1.XA4.LCK_N AVSS 1.25521f
C4499 XA2.XA1.XA5.MN2.S AVSS 0.049396f
C4500 XA1.XA1.XA5.MN2.S AVSS 0.049396f
C4501 XA0.XA1.XA5.MN1.S AVSS 0.10078f
C4502 XA0.XA1.XA4.LCK_N AVSS 1.2666f
C4503 XA0.XA1.XA5.MN2.S AVSS 0.049396f
C4504 a_19982_42588# AVSS 0.4015f $ **FLOATING
C4505 a_18614_42588# AVSS 0.40162f $ **FLOATING
C4506 a_14942_42588# AVSS 0.40162f $ **FLOATING
C4507 a_13574_42588# AVSS 0.40162f $ **FLOATING
C4508 a_9902_42588# AVSS 0.401051f $ **FLOATING
C4509 a_8534_42588# AVSS 0.399959f $ **FLOATING
C4510 a_4862_42588# AVSS 0.400568f $ **FLOATING
C4511 a_3494_42588# AVSS 0.399691f $ **FLOATING
C4512 a_n178_42588# AVSS 0.401905f $ **FLOATING
C4513 XA0.CMP_OP AVSS 16.905f
C4514 a_23654_43116# AVSS 0.425494f $ **FLOATING
C4515 XA8.XA2.A AVSS 2.24226f
C4516 XA7.XA2.A AVSS 2.22341f
C4517 XA6.XA2.A AVSS 2.22305f
C4518 XA5.XA2.A AVSS 2.22341f
C4519 XA4.XA2.A AVSS 2.2181f
C4520 XA3.XA2.A AVSS 2.20215f
C4521 XA2.XA2.A AVSS 2.21221f
C4522 XA1.XA2.A AVSS 2.19894f
C4523 XA0.XA2.A AVSS 2.22411f
C4524 a_19982_43468# AVSS 0.426697f $ **FLOATING
C4525 a_18614_43468# AVSS 0.426697f $ **FLOATING
C4526 a_14942_43468# AVSS 0.426697f $ **FLOATING
C4527 a_13574_43468# AVSS 0.426697f $ **FLOATING
C4528 a_9902_43468# AVSS 0.426128f $ **FLOATING
C4529 a_8534_43468# AVSS 0.425036f $ **FLOATING
C4530 a_4862_43468# AVSS 0.425644f $ **FLOATING
C4531 a_3494_43468# AVSS 0.424768f $ **FLOATING
C4532 a_n178_43468# AVSS 0.426982f $ **FLOATING
C4533 XA0.CMP_ON AVSS 20.8286f
C4534 a_23654_43996# AVSS 0.42719f $ **FLOATING
C4535 XA8.CN1 AVSS 3.01685f
C4536 XA7.CN1 AVSS 2.99708f
C4537 XA6.CN1 AVSS 2.99623f
C4538 XA5.CN1 AVSS 2.99708f
C4539 XA4.CN1 AVSS 2.99599f
C4540 XA3.CN1 AVSS 9.974581f
C4541 XA2.CN1 AVSS 10.5726f
C4542 XA1.CN1 AVSS 9.95499f
C4543 a_19982_44348# AVSS 0.427289f $ **FLOATING
C4544 a_18614_44348# AVSS 0.427289f $ **FLOATING
C4545 a_14942_44348# AVSS 0.427289f $ **FLOATING
C4546 a_13574_44348# AVSS 0.427289f $ **FLOATING
C4547 a_9902_44348# AVSS 0.427289f $ **FLOATING
C4548 a_8534_44348# AVSS 0.427289f $ **FLOATING
C4549 a_4862_44348# AVSS 0.427289f $ **FLOATING
C4550 a_3494_44348# AVSS 0.427289f $ **FLOATING
C4551 a_n178_44348# AVSS 0.428057f $ **FLOATING
C4552 XA20.XA2.N1 AVSS 1.61009f
C4553 XA20.XA3.N2 AVSS 0.331373f
C4554 XA8.XA1.CHL_OP AVSS 3.27318f
C4555 XA7.XA1.CHL_OP AVSS 3.24106f
C4556 XA6.XA1.CHL_OP AVSS 3.24233f
C4557 XA5.XA1.CHL_OP AVSS 3.24106f
C4558 XA4.XA1.CHL_OP AVSS 3.23938f
C4559 XA3.XA1.CHL_OP AVSS 3.23799f
C4560 XA2.XA1.CHL_OP AVSS 3.2392f
C4561 XA1.XA1.CHL_OP AVSS 3.23799f
C4562 XA0.XA1.CHL_OP AVSS 3.3272f
C4563 XA20.XA2.VMR AVSS 2.70278f
C4564 XA20.XA2.CO AVSS 2.70435f
C4565 a_19982_45228# AVSS 0.426697f $ **FLOATING
C4566 a_18614_45228# AVSS 0.426697f $ **FLOATING
C4567 a_14942_45228# AVSS 0.426697f $ **FLOATING
C4568 a_13574_45228# AVSS 0.426697f $ **FLOATING
C4569 a_9902_45228# AVSS 0.426697f $ **FLOATING
C4570 a_8534_45228# AVSS 0.426697f $ **FLOATING
C4571 a_4862_45228# AVSS 0.426697f $ **FLOATING
C4572 a_3494_45228# AVSS 0.426697f $ **FLOATING
C4573 a_n178_45228# AVSS 0.4277f $ **FLOATING
C4574 a_23654_45404# AVSS 0.404684f $ **FLOATING
C4575 XA8.CP0 AVSS 3.07901f
C4576 XA7.CP0 AVSS 3.07648f
C4577 XA6.CP0 AVSS 3.07638f
C4578 XA5.CP0 AVSS 3.07648f
C4579 XA4.CP0 AVSS 3.07638f
C4580 XA3.CP0 AVSS 6.31197f
C4581 XA2.CP0 AVSS 6.44611f
C4582 XA1.CP0 AVSS 12.127901f
C4583 XA0.CP0 AVSS 16.1686f
C4584 a_19982_46108# AVSS 0.427411f $ **FLOATING
C4585 a_18614_46108# AVSS 0.427356f $ **FLOATING
C4586 a_14942_46108# AVSS 0.427356f $ **FLOATING
C4587 a_13574_46108# AVSS 0.427356f $ **FLOATING
C4588 a_9902_46108# AVSS 0.427356f $ **FLOATING
C4589 a_8534_46108# AVSS 0.427356f $ **FLOATING
C4590 a_4862_46108# AVSS 0.427356f $ **FLOATING
C4591 a_3494_46108# AVSS 0.427356f $ **FLOATING
C4592 a_n178_46108# AVSS 0.428328f $ **FLOATING
C4593 XA20.XA4.MP0.S AVSS 0.545672f
C4594 XA8.XA6.MN1.S AVSS 0.168832f
C4595 XA8.CN0 AVSS 0.70463f
C4596 XA7.XA6.MN1.S AVSS 0.150197f
C4597 a_23654_46812# AVSS 0.395265f $ **FLOATING
C4598 XA7.CN0 AVSS 8.63576f
C4599 XA6.XA6.MN1.S AVSS 0.150197f
C4600 XA6.CN0 AVSS 6.24771f
C4601 XA8.XA6.MN3.S AVSS 0.094305f
C4602 XA7.XA6.MN3.S AVSS 0.102759f
C4603 XA5.XA6.MN1.S AVSS 0.150197f
C4604 XA5.CN0 AVSS 4.94098f
C4605 XA4.XA6.MN1.S AVSS 0.150197f
C4606 XA4.CN0 AVSS 6.34921f
C4607 XA6.XA6.MN3.S AVSS 0.102759f
C4608 XA5.XA6.MN3.S AVSS 0.102759f
C4609 XA3.XA6.MN1.S AVSS 0.150197f
C4610 XA3.CN0 AVSS 4.51265f
C4611 XA2.XA6.MN1.S AVSS 0.150197f
C4612 XA2.CN0 AVSS 4.83638f
C4613 XA4.XA6.MN3.S AVSS 0.102759f
C4614 XA3.XA6.MN3.S AVSS 0.102759f
C4615 XA1.XA6.MN1.S AVSS 0.150197f
C4616 XA1.CN0 AVSS 10.6047f
C4617 XA0.XA6.MN1.S AVSS 0.150572f
C4618 XA0.CN0 AVSS 14.822598f
C4619 XA2.XA6.MN3.S AVSS 0.102759f
C4620 XA1.XA6.MN3.S AVSS 0.102759f
C4621 XA0.XA6.MN3.S AVSS 0.103205f
C4622 XA0.CP1 AVSS 14.794499f
C4623 a_19982_46988# AVSS 0.393747f $ **FLOATING
C4624 a_18614_46988# AVSS 0.395238f $ **FLOATING
C4625 a_14942_46988# AVSS 0.395238f $ **FLOATING
C4626 a_13574_46988# AVSS 0.395238f $ **FLOATING
C4627 a_9902_46988# AVSS 0.395238f $ **FLOATING
C4628 a_8534_46988# AVSS 0.395238f $ **FLOATING
C4629 a_4862_46988# AVSS 0.395238f $ **FLOATING
C4630 a_3494_46988# AVSS 0.395238f $ **FLOATING
C4631 a_n178_46988# AVSS 0.396006f $ **FLOATING
C4632 XA20.XA1.CK AVSS 4.76072f
C4633 a_23654_47164# AVSS 0.395827f $ **FLOATING
C4634 XA8.ENO AVSS 1.79727f
C4635 XA7.ENO AVSS 4.52797f
C4636 XA6.ENO AVSS 4.34408f
C4637 XA5.ENO AVSS 4.47264f
C4638 XA4.ENO AVSS 4.35438f
C4639 XA4.EN AVSS 4.49527f
C4640 XA2.ENO AVSS 4.40632f
C4641 XA1.ENO AVSS 4.4603f
C4642 XA0.ENO AVSS 4.40615f
C4643 XA20.XA10.MN1.S AVSS 0.097455f
C4644 a_19982_47340# AVSS 0.389919f $ **FLOATING
C4645 a_18614_47340# AVSS 0.389919f $ **FLOATING
C4646 a_14942_47340# AVSS 0.389919f $ **FLOATING
C4647 a_13574_47340# AVSS 0.389919f $ **FLOATING
C4648 a_9902_47340# AVSS 0.389919f $ **FLOATING
C4649 a_8534_47340# AVSS 0.389919f $ **FLOATING
C4650 a_4862_47340# AVSS 0.389919f $ **FLOATING
C4651 a_3494_47340# AVSS 0.389919f $ **FLOATING
C4652 a_n178_47340# AVSS 0.390688f $ **FLOATING
C4653 XA20.XA1.CKN AVSS 5.03067f
C4654 XA7.DONE AVSS 0.236186f
C4655 XA6.DONE AVSS 0.236186f
C4656 XA5.DONE AVSS 0.236186f
C4657 XA4.DONE AVSS 0.236186f
C4658 XA3.DONE AVSS 0.236186f
C4659 XA2.DONE AVSS 0.236186f
C4660 XA1.DONE AVSS 0.236186f
C4661 XA0.DONE AVSS 0.236186f
C4662 a_23654_47692# AVSS 0.397011f $ **FLOATING
C4663 a_19982_47692# AVSS 0.391328f $ **FLOATING
C4664 a_18614_47692# AVSS 0.393098f $ **FLOATING
C4665 a_14942_47692# AVSS 0.393098f $ **FLOATING
C4666 a_13574_47692# AVSS 0.393098f $ **FLOATING
C4667 a_9902_47692# AVSS 0.393098f $ **FLOATING
C4668 a_8534_47692# AVSS 0.393098f $ **FLOATING
C4669 a_4862_47692# AVSS 0.393098f $ **FLOATING
C4670 a_3494_47692# AVSS 0.393098f $ **FLOATING
C4671 a_n178_47692# AVSS 0.393899f $ **FLOATING
C4672 XA8.XA8.A AVSS 1.5261f
C4673 XA8.XA9.MN1.S AVSS 0.113648f
C4674 XA20.XA10.A AVSS 1.07576f
C4675 XA8.XA6.Y AVSS 1.56237f
C4676 XA7.XA9.MN1.S AVSS 0.113648f
C4677 XA7.XA8.A AVSS 1.52787f
C4678 XA7.XA6.Y AVSS 1.56895f
C4679 XA6.XA8.A AVSS 1.52787f
C4680 XA6.XA9.MN1.S AVSS 0.113648f
C4681 XA6.XA6.Y AVSS 1.57794f
C4682 XA5.XA9.MN1.S AVSS 0.113648f
C4683 XA5.XA8.A AVSS 1.52787f
C4684 XA5.XA6.Y AVSS 1.56895f
C4685 XA4.XA8.A AVSS 1.52787f
C4686 XA4.XA9.MN1.S AVSS 0.113648f
C4687 XA4.XA6.Y AVSS 1.57794f
C4688 XA3.XA9.MN1.S AVSS 0.113648f
C4689 XA3.XA8.A AVSS 1.52787f
C4690 XA3.XA6.Y AVSS 1.56895f
C4691 XA2.XA8.A AVSS 1.52787f
C4692 XA2.XA9.MN1.S AVSS 0.113648f
C4693 XA2.XA6.Y AVSS 1.57794f
C4694 XA1.XA9.MN1.S AVSS 0.113648f
C4695 XA1.XA8.A AVSS 1.52787f
C4696 XA1.XA6.Y AVSS 1.56895f
C4697 XA0.XA8.A AVSS 1.53082f
C4698 XA0.XA9.MN1.S AVSS 0.113648f
C4699 XA0.XA6.Y AVSS 1.62644f
C4700 a_23654_48220# AVSS 0.416084f $ **FLOATING
C4701 a_19982_48220# AVSS 0.391706f $ **FLOATING
C4702 a_18614_48220# AVSS 0.391706f $ **FLOATING
C4703 a_14942_48220# AVSS 0.391706f $ **FLOATING
C4704 a_13574_48220# AVSS 0.391706f $ **FLOATING
C4705 a_9902_48220# AVSS 0.391706f $ **FLOATING
C4706 a_8534_48220# AVSS 0.391706f $ **FLOATING
C4707 a_4862_48220# AVSS 0.391706f $ **FLOATING
C4708 a_3494_48220# AVSS 0.391706f $ **FLOATING
C4709 a_n178_48220# AVSS 0.392709f $ **FLOATING
C4710 XA20.XA10.B AVSS 0.792299f
C4711 XA8.XA10.A AVSS 0.898521f
C4712 XA7.XA10.A AVSS 0.898521f
C4713 XA6.XA10.A AVSS 0.898521f
C4714 XA5.XA10.A AVSS 0.898521f
C4715 XA4.XA10.A AVSS 0.898521f
C4716 XA3.XA10.A AVSS 0.898521f
C4717 XA2.XA10.A AVSS 0.898521f
C4718 XA1.XA10.A AVSS 0.898521f
C4719 XA0.XA10.A AVSS 0.899973f
C4720 a_23654_48572# AVSS 0.476259f $ **FLOATING
C4721 a_19982_48572# AVSS 0.395129f $ **FLOATING
C4722 a_18614_48572# AVSS 0.394787f $ **FLOATING
C4723 a_14942_48572# AVSS 0.395129f $ **FLOATING
C4724 a_13574_48572# AVSS 0.394787f $ **FLOATING
C4725 a_9902_48572# AVSS 0.395129f $ **FLOATING
C4726 a_8534_48572# AVSS 0.394787f $ **FLOATING
C4727 a_4862_48572# AVSS 0.395129f $ **FLOATING
C4728 a_3494_48572# AVSS 0.394787f $ **FLOATING
C4729 a_n178_48572# AVSS 0.396133f $ **FLOATING
C4730 a_23654_48924# AVSS 0.542949f $ **FLOATING
C4731 a_22502_48924# AVSS 0.090319f $ **FLOATING
C4732 XA8.XA10.Y AVSS 0.894759f
C4733 XA7.XA10.Y AVSS 0.886801f
C4734 XA6.XA10.Y AVSS 0.894775f
C4735 XA5.XA10.Y AVSS 0.886801f
C4736 XA4.XA10.Y AVSS 0.894775f
C4737 XA3.XA10.Y AVSS 0.886801f
C4738 XA2.XA10.Y AVSS 0.894775f
C4739 XA1.XA10.Y AVSS 0.886801f
C4740 XA0.XA10.Y AVSS 0.896291f
C4741 XB1.TIE_L AVSS 35.6477f
C4742 a_19982_49100# AVSS 0.413874f $ **FLOATING
C4743 a_18614_49100# AVSS 0.413588f $ **FLOATING
C4744 a_14942_49100# AVSS 0.413874f $ **FLOATING
C4745 a_13574_49100# AVSS 0.413588f $ **FLOATING
C4746 a_9902_49100# AVSS 0.413874f $ **FLOATING
C4747 a_8534_49100# AVSS 0.413588f $ **FLOATING
C4748 a_4862_49100# AVSS 0.413874f $ **FLOATING
C4749 a_3494_49100# AVSS 0.413588f $ **FLOATING
C4750 a_n178_49100# AVSS 0.414878f $ **FLOATING
C4751 XA8.XA11.Y AVSS 1.12045f
C4752 XA8.CEO AVSS 1.22181f
C4753 XA7.XA11.Y AVSS 1.07541f
C4754 XA7.CEO AVSS 1.73212f
C4755 XA6.XA11.Y AVSS 1.11767f
C4756 XA6.CEO AVSS 1.55142f
C4757 XA5.XA11.Y AVSS 1.07541f
C4758 XA5.CEO AVSS 1.73122f
C4759 XA4.XA11.Y AVSS 1.11767f
C4760 XA4.CEO AVSS 1.55142f
C4761 XA3.XA11.Y AVSS 1.07541f
C4762 XA4.CEIN AVSS 1.73122f
C4763 XA2.XA11.Y AVSS 1.11767f
C4764 XA2.CEO AVSS 1.55142f
C4765 XA1.XA11.Y AVSS 1.07541f
C4766 XA1.CEO AVSS 1.73122f
C4767 XA0.XA11.Y AVSS 1.11905f
C4768 XA0.CEO AVSS 1.54913f
C4769 a_19982_49452# AVSS 0.474508f $ **FLOATING
C4770 a_18614_49452# AVSS 0.476112f $ **FLOATING
C4771 a_14942_49452# AVSS 0.474508f $ **FLOATING
C4772 a_13574_49452# AVSS 0.476112f $ **FLOATING
C4773 a_9902_49452# AVSS 0.474508f $ **FLOATING
C4774 a_8534_49452# AVSS 0.476112f $ **FLOATING
C4775 a_4862_49452# AVSS 0.474508f $ **FLOATING
C4776 a_3494_49452# AVSS 0.476112f $ **FLOATING
C4777 a_n178_49452# AVSS 0.47548f $ **FLOATING
C4778 a_21134_49804# AVSS 0.097214f $ **FLOATING
C4779 a_19982_49804# AVSS 0.546762f $ **FLOATING
C4780 a_18614_49804# AVSS 0.545607f $ **FLOATING
C4781 a_17462_49804# AVSS 0.096044f $ **FLOATING
C4782 a_16094_49804# AVSS 0.096044f $ **FLOATING
C4783 a_14942_49804# AVSS 0.546762f $ **FLOATING
C4784 a_13574_49804# AVSS 0.545607f $ **FLOATING
C4785 a_12422_49804# AVSS 0.096044f $ **FLOATING
C4786 a_11054_49804# AVSS 0.096044f $ **FLOATING
C4787 a_9902_49804# AVSS 0.546762f $ **FLOATING
C4788 a_8534_49804# AVSS 0.545607f $ **FLOATING
C4789 a_7382_49804# AVSS 0.096044f $ **FLOATING
C4790 a_6014_49804# AVSS 0.096044f $ **FLOATING
C4791 a_4862_49804# AVSS 0.546762f $ **FLOATING
C4792 a_3494_49804# AVSS 0.545607f $ **FLOATING
C4793 a_2342_49804# AVSS 0.096044f $ **FLOATING
C4794 a_974_49804# AVSS 0.096044f $ **FLOATING
C4795 a_n178_49804# AVSS 0.547733f $ **FLOATING
.ends

