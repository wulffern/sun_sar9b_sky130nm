magic
tech sky130A
magscale 1 2
timestamp 1708902000
<< checkpaint >>
rect 0 0 184 68
<< m2 >>
rect 0 0 184 68
<< v2 >>
rect 12 6 68 62
rect 116 6 172 62
<< m3 >>
rect 0 0 184 68
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 184 68
<< end >>
