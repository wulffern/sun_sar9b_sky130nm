magic
tech sky130A
timestamp 1708968222
<< locali >>
rect 84 1562 720 1596
rect 84 1332 118 1562
rect 314 1347 432 1381
rect 0 1298 118 1332
rect 199 775 233 1337
rect 314 1205 348 1347
rect 378 1259 550 1293
rect 314 1171 432 1205
rect 314 1029 348 1171
rect 516 1117 550 1259
rect 432 1083 550 1117
rect 314 995 432 1029
rect 314 853 348 995
rect 516 941 550 1083
rect 432 907 550 941
rect 314 819 432 853
rect 314 677 348 819
rect 516 765 550 907
rect 432 731 550 765
rect 314 643 432 677
rect 199 71 233 633
rect 314 501 348 643
rect 378 555 550 589
rect 314 467 432 501
rect 314 325 348 467
rect 516 413 550 555
rect 1710 423 1818 457
rect 432 379 550 413
rect 314 291 432 325
rect 314 149 348 291
rect 516 237 550 379
rect 882 247 990 281
rect 432 203 550 237
rect 314 115 432 149
rect 516 61 550 203
rect 432 27 550 61
<< metal1 >>
rect 300 1435 1152 1469
rect 300 1337 334 1435
rect 216 1303 334 1337
rect 1020 1100 1548 1134
rect 1020 897 1054 1100
rect 936 863 1054 897
rect 1494 819 1710 853
rect 516 643 1152 677
rect 516 501 550 643
rect 432 467 550 501
rect 1632 423 1764 457
rect 1632 325 1666 423
rect 1548 291 1666 325
<< metal2 >>
rect 716 907 1152 941
rect 716 457 750 907
rect 936 775 1054 809
rect 216 423 750 457
rect 1020 342 1054 775
rect 1548 555 1666 589
rect 1020 308 1152 342
rect 1632 14 1666 555
rect 1632 -20 2188 14
<< metal3 >>
rect 838 1435 930 1469
rect 394 115 486 149
rect 1098 0 1190 2400
rect 1494 0 1586 2400
rect 2078 1340 3924 1374
rect 2078 853 2112 1340
rect 1756 819 2112 853
use SUNSAR_NCHDLR  M1
timestamp 1708902000
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_NCHDLR  M2
timestamp 1708902000
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNSAR_NCHDLR  M3
timestamp 1708902000
transform 1 0 0 0 1 352
box -90 -66 630 242
use SUNSAR_NCHDLR  M4
timestamp 1708902000
transform 1 0 0 0 1 528
box -90 -66 630 242
use SUNSAR_NCHDLR  M5
timestamp 1708902000
transform 1 0 0 0 1 704
box -90 -66 630 242
use SUNSAR_NCHDLR  M6
timestamp 1708902000
transform 1 0 0 0 1 880
box -90 -66 630 242
use SUNSAR_NCHDLR  M7
timestamp 1708902000
transform 1 0 0 0 1 1056
box -90 -66 630 242
use SUNSAR_NCHDLR  M8
timestamp 1708902000
transform 1 0 0 0 1 1232
box -90 -66 630 242
use SUNSAR_IVX1_CV  XA0
timestamp 1708968222
transform 1 0 720 0 1 176
box -90 -66 1350 242
use SUNSAR_TIEH_CV  XA1
timestamp 1708968222
transform 1 0 720 0 1 968
box -90 -66 1350 242
use SUNSAR_TIEL_CV  XA2
timestamp 1708968222
transform 1 0 720 0 1 1320
box -90 -66 1350 242
use SUNSAR_TGPD_CV  XA3
timestamp 1708968222
transform 1 0 720 0 1 352
box -90 -66 1350 418
use SUNSAR_SARBSSWCTRL_CV  XA4
timestamp 1708968222
transform 1 0 720 0 1 704
box -90 -66 1350 330
use SUNSAR_TAPCELLB_CV  XA5
timestamp 1708968222
transform 1 0 720 0 1 1496
box -90 -66 1350 242
use SUNSAR_TAPCELLB_CV  XA5b
timestamp 1708968222
transform 1 0 720 0 1 0
box -90 -66 1350 242
use SUNSAR_TAPCELLB_CV  XA7
timestamp 1708968222
transform 1 0 720 0 1 1144
box -90 -66 1350 242
use SUNSAR_CAP_BSSW5_CV  XCAPB1
timestamp 1708968222
transform 1 0 2088 0 1 0
box -10 -20 3682 2340
use SUNSAR_cut_M1M2_2x1  xcut0
timestamp 1708902000
transform 1 0 1494 0 1 819
box 0 0 92 34
use SUNSAR_cut_M2M4_2x1  xcut1
timestamp 1708902000
transform 1 0 1710 0 1 819
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut2
timestamp 1708902000
transform 1 0 1494 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut3
timestamp 1708902000
transform 1 0 1710 0 1 423
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut4
timestamp 1708902000
transform 1 0 882 0 1 775
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut5
timestamp 1708902000
transform 1 0 1098 0 1 308
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut6
timestamp 1708902000
transform 1 0 162 0 1 1303
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut7
timestamp 1708902000
transform 1 0 1098 0 1 1435
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut8
timestamp 1708902000
transform 1 0 882 0 1 863
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut9
timestamp 1708902000
transform 1 0 1494 0 1 1100
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut10
timestamp 1708902000
transform 1 0 378 0 1 467
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut11
timestamp 1708902000
transform 1 0 1098 0 1 643
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut12
timestamp 1708902000
transform 1 0 1114 0 1 907
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut13
timestamp 1708902000
transform 1 0 178 0 1 423
box 0 0 92 34
use SUNSAR_cut_M1M3_2x1  xcut14
timestamp 1708902000
transform 1 0 1494 0 1 555
box 0 0 92 34
use SUNSAR_cut_M3M4_2x1  xcut15
timestamp 1708902000
transform 1 0 2142 0 1 -20
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut16
timestamp 1708902000
transform 1 0 394 0 1 115
box 0 0 92 34
use SUNSAR_cut_M2M4_2x1  xcut17
timestamp 1708902000
transform 1 0 838 0 1 1435
box 0 0 92 34
<< labels >>
flabel metal3 s 394 115 486 149 0 FreeSans 200 0 0 0 VI
port 1 nsew signal bidirectional
flabel metal3 s 838 1435 930 1469 0 FreeSans 200 0 0 0 TIE_L
port 4 nsew signal bidirectional
flabel locali s 882 247 990 281 0 FreeSans 200 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 1710 423 1818 457 0 FreeSans 200 0 0 0 CKN
port 3 nsew signal bidirectional
flabel locali s 378 555 486 589 0 FreeSans 200 0 0 0 VO1
port 5 nsew signal bidirectional
flabel locali s 378 1259 486 1293 0 FreeSans 200 0 0 0 VO2
port 6 nsew signal bidirectional
flabel metal3 s 1494 0 1586 2400 0 FreeSans 200 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel metal3 s 1098 0 1190 2400 0 FreeSans 200 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 5724 2400
<< end >>
