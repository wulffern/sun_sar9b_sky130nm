**********************************************************************
**        Copyright (c) 2016 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2016-11-16
** *******************************************************************


.subckt TIEH_CV Y BULKP BULKN AVDD AVSS
MN0 A A AVSS BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
.ends

.subckt TIEL_CV Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MP0 A A AVDD BULKP PCHDL
.ends TIEL_CV


.subckt IVX1_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
.ends

.subckt TIVX1_CV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
.ends

.subckt IVX2_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
.ends

.subckt IVX4_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
MP2 Y A AVDD BULKP PCHDL
MP3 AVDD A Y BULKP PCHDL
.ends IVX4_CV

.subckt IVX8_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MN4 Y A AVSS BULKN NCHDL
MN5 AVSS A Y BULKN NCHDL
MN6 Y A AVSS BULKN NCHDL
MN7 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
MP2 Y A AVDD BULKP PCHDL
MP3 AVDD A Y BULKP PCHDL
MP4 Y A AVDD BULKP PCHDL
MP5 AVDD A Y BULKP PCHDL
MP6 Y A AVDD BULKP PCHDL
MP7 AVDD A Y BULKP PCHDL
.ends IVX8_CV

.subckt BFX1_CV A Y BULKP BULKN AVDD AVSS
MN0 AVSS A B BULKN NCHDL
MN1 Y B AVSS BULKN NCHDL
MP0 AVDD A B BULKP PCHDL
MP1 Y B AVDD BULKP PCHDL
.ends BFX1_CV





*-----------------------------------------------------------------------------
* NAND/NOR
*-----------------------------------------------------------------------------

.subckt NRX1_CV A B Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN  NCHDL
MN1 AVSS B Y BULKN  NCHDL
MP0 N1 A AVDD BULKP PCHDL
MP1 Y B N1 BULKP PCHDL
.ends NRX1_CV

.subckt NDX1_CV A B Y BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN NCHDL
MN1 Y B N1 BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD B Y BULKP PCHDL
.ends NDX1_CV

.subckt ORX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS  NRX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS  IVX1_CV
.ends

.subckt ANX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS IVX1_CV
.ends


.subckt IVTRIX1_CV A C CN Y  BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN NCHDL
MN1 Y C N1 BULKN NCHDL
MP0 N2 A AVDD BULKP PCHDL
MP1 Y CN N2 BULKP PCHDL
.ends IVTRIX1_CV

.subckt NDTRIX1_CV A C CN RN Y BULKP BULKN AVDD AVSS
MN2 N1 RN AVSS BULKN NCHDL
MN0 N2 A N1 BULKN NCHDL
MN1 Y C N2 BULKN NCHDL
MP2 AVDD RN N2 BULKP PCHDL
MP0 N2 A AVDD BULKP PCHDL
MP1 Y CN N2 BULKP PCHDL
.ends


.subckt DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS AVDD AVSS NDX1_CV
XA2 CKN CKB AVDD AVSS AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS AVDD AVSS IVTRIX1_CV
XA5 A0 A1 AVDD AVSS AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS AVDD AVSS NDTRIX1_CV
XA8 QN Q AVDD AVSS AVDD AVSS IVX1_CV

.ends


.SUBCKT SCX1_CV A Y BULKP BULKN  AVDD AVSS
XA2 N1 A AVSS BULKN  NCHDL
XA3 SCO A N1 BULKN  NCHDL
XA4a AVDD SCO N1 BULKN  NCHDL
XA4b AVDD SCO N1 BULKN  NCHDL
XA5 Y SCO AVSS BULKN  NCHDL

XB0 N2 A AVDD BULKP  PCHDL
XB1 SCO A N2 BULKP  PCHDL
XB3a N2 SCO AVSS BULKP  PCHDL
XB3b N2 SCO AVSS BULKP  PCHDL
XB4 Y SCO AVDD AVSS  PCHDL
.ends


*-----------------------------------------------------------------------------
* SAR unit logic cells
*---------------------------------------------------------------------------




.subckt DMY_CV
MN0  NCHDLDMY
MP0  PCHDLDMY
.ends DNY_CV


.SUBCKT TAPCELLB_CV AVDD AVSS
MN1 AVSS AVSS AVSS AVSS  NCHDL
MP1 AVDD AVDD AVDD AVDD  PCHDL
.ENDS


.subckt SWX2_CV A Y VREF AVSS BULKP BULKN
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MP0 Y A VREF BULKP PCHDL
MP1 VREF A Y BULKP PCHDL
.ends SWX2_CV


.subckt SWX4_CV A Y VREF AVSS BULKP BULKN
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MP0 Y A VREF BULKP PCHDL
MP1 VREF A Y BULKP PCHDL
MP2 Y A VREF BULKP PCHDL
MP3 VREF A Y BULKP PCHDL
.ends IVX4_CV

.subckt TGPD_CV C A B BULKP BULKN AVDD AVSS
MN0 AVSS C CN BULKN NCHDL
MN1 B C AVSS BULKN NCHDL
MN2 A CN B BULKN NCHDL
MP0 AVDD C CN BULKP PCHDL
MP1_DMY B AVDD AVDD BULKP PCHDL
MP2 A C B BULKP PCHDL
.ends


.subckt SARBSSWCTRL_CV C GN GNG TIE_H  BULKP BULKN AVDD AVSS
MN0 N1 C AVSS BULKN NCHDL
MN1 GN TIE_H N1 BULKN NCHDL
MP0 GNG C GN BULKP PCHDL
MP1 AVDD GN GNG BULKP PCHDL
.ends

.SUBCKT SAREMX1_CV A  B EN ENO RST_N BULKP BULKN AVDD AVSS
MN0 N3 EN AM BULKN  NCHDL
MN1 N3 B AVSS BULKN  NCHDL
MN2 AVSS A N3 BULKN  NCHDL
MN3 ENO AM AVSS BULKN  NCHDL
MP0 AVDD RST_N AM BULKP PCHDL
MP1 N2 B ENO BULKP  PCHDL
MP2 N1 A N2 BULKP  PCHDL
MP3 AVDD AM N1 BULKP  PCHDL
.ENDS

.SUBCKT SARLTX1_CV A CHL RST_N EN LCK_N BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN  NCHDL
MN1 N3 LCK_N N1 BULKN  NCHDL
MN2 CHL EN N3 BULKN  NCHDL
MP0 NP2 RST_N AVDD BULKP PCHDL
MP1 NP1 RST_N NP2 BULKP PCHDL
MP2 CHL RST_N NP1 BULKP PCHDL
.ENDS

.SUBCKT SARCEX1_CV A B Y RST  BULKP BULKN AVDD AVSS
MN0 N4 RST AVSS BULKN  NCHDL
MN1 AVSS RST N4 BULKN  NCHDL
MN2 N1 RST AVSS BULKN  NCHDL
MN3 Y RST N1 BULKN  NCHDL

MP0 N2 A Y BULKP PCHDL
MP1 AVDD A N2 BULKP PCHDL
MP2 N3 B AVDD BULKP PCHDL
MP3 Y B N3 BULKP PCHDL
.ENDS

.SUBCKT SARCMPHX1_CV CI CK CO VMR N1 N2 BULKP BULKN AVDD AVSS
MN0  N1 CK AVSS BULKN NCHDL
MN1  N2 CI N1   BULKN NCHDL
MN2  N1 CI N2   BULKN NCHDL
MN3  N2 CI N1   BULKN NCHDL
MN4  N1 CI N2   BULKN NCHDL
MN5  N2 CI N1   BULKN NCHDL
MN6  CO VMR N2   BULKN NCHDL

MP0  AVDD CK N1 BULKP PCHDL
MP1  N2 CK AVDD BULKP PCHDL
MP2  AVDD AVDD N2 BULKP PCHDL
MP3  CO CK AVDD BULKP PCHDL
MP4  AVDD VMR CO BULKP PCHDL
MP5  CO VMR AVDD BULKP PCHDL
MP6  AVDD VMR CO BULKP PCHDL
.ENDS SARCMPHX1_CV


.SUBCKT SARKICKHX1_CV CI CK CKN BULKP BULKN AVDD AVSS
MN0  N1 CKN AVSS BULKN NCHDL
MN1  N1 CI N1   BULKN NCHDL
MN2  N1 CI N1   BULKN NCHDL
MN3  N1 CI N1   BULKN NCHDL
MN4  N1 CI N1   BULKN NCHDL
MN5  N1 CI N1   BULKN NCHDL
MN6  AVDD CK N1   BULKN NCHDL

MP0  AVDD CKN N1 BULKP PCHDL
MP1_DMY AVDD AVDD AVDD BULKP PCHDL
MP2_DMY AVDD AVDD AVDD BULKP PCHDL
MP3_DMY AVDD AVDD AVDD BULKP PCHDL
MP4_DMY AVDD AVDD AVDD BULKP PCHDL
MP5_DMY AVDD AVDD AVDD BULKP PCHDL
MP6_DMY  AVDD AVDD AVDD BULKP PCHDL
.ENDS SARKICKHX1_CV


*-----------------------------------------------------------------------------
* SAR composite logic cells
*---------------------------------------------------------------------------

.subckt TEST_CV A Y AVDD AVSS
XA5 AVDD AVSS TAPCELLB_CV
XA2 A Y AVDD AVSS TIVX1_CV
.ends


.SUBCKT CAP_BSSW5_CV A B
XCAPB A B CAP_BSSW_CV M=5
.ENDS

.SUBCKT SARBSSW_CV VI CK CKN TIE_L VO1 VO2 AVDD AVSS

M1 VI GN VO1 AVSS NCHDLR
M2 VI GN VO1 AVSS NCHDLR
M3 VI GN VO1 AVSS NCHDLR
M4 VI GN VO1 AVSS NCHDLR
M5 VI TIE_L VO2 AVSS NCHDLR
M6 VI TIE_L VO2 AVSS NCHDLR
M7 VI TIE_L VO2 AVSS NCHDLR
M8 VI TIE_L VO2 AVSS NCHDLR

XA5b AVDD AVSS TAPCELLB_CV
XA0 CK CKN AVDD AVSS AVDD AVSS IVX1_CV
XA3 CKN VI VS AVDD AVSS AVDD AVSS TGPD_CV
XA4 CKN GN GNG TIE_H AVDD AVSS AVDD AVSS SARBSSWCTRL_CV
XA1 TIE_H AVDD AVSS AVDD AVSS TIEH_CV
XA7 AVDD AVSS TAPCELLB_CV
XA2 TIE_L AVDD AVSS AVDD AVSS TIEL_CV
XA5 AVDD AVSS TAPCELLB_CV


XCAPB1 GNG VS CAP_BSSW5_CV xoffset=3
*XCAPB2 GNG VS CAP_BSSW_CV M=4
*XCAP GNG VS CAPX10_CV
*XCAPB GNG VS CAPX1_CV M=7
*XCAPC GNG VS CAPX1_CV M=7

.ENDS

.SUBCKT SARCMPX1_CV CPI CNI CPO CNO CK_CMP CK_SAMPLE DONE AVDD AVSS
*XA0a DMY_CV
XA0 AVDD AVSS TAPCELLB_CV
XA1 CPI CK_B CK_N AVDD AVSS AVDD AVSS SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS AVDD AVSS SARCMPHX1_CV
XA2a CPO_I CPO AVDD AVSS AVDD AVSS IVX4_CV
XA3a CNO_I CNO AVDD AVSS AVDD AVSS IVX4_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS  AVDD AVSS SARCMPHX1_CV
XA4 CNI CK_B CK_N AVDD AVSS AVDD AVSS SARKICKHX1_CV
XA9 CK_N CK_B AVDD AVSS AVDD AVSS IVX1_CV
XA10 DONE_N CK_A CK_N AVDD AVSS AVDD AVSS NDX1_CV
XA11 CK_SAMPLE DONE DONE_N AVDD AVSS AVDD AVSS NRX1_CV
XA12 CK_CMP CK_A AVDD AVSS AVDD AVSS IVX1_CV
XA13 AVDD AVSS TAPCELLB_CV
*XA14 DMY_CV
.ENDS

.SUBCKT SARCMPX2_CV CPI CNI CPO CNO CK_CMP CK_SAMPLE DONE AVDD AVSS
*XA0a DMY_CV
XA0 AVDD AVSS TAPCELLB_CV
XA1 CPI CK_B CK_N AVDD AVSS AVDD AVSS SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS AVDD AVSS SARCMPHX1_CV
XA2a CPO_I CPO AVDD AVSS AVDD AVSS IVX2_CV
XA3a CNO_I CNO AVDD AVSS AVDD AVSS IVX2_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS  AVDD AVSS SARCMPHX1_CV
XA4 CNI CK_B CK_N AVDD AVSS AVDD AVSS SARKICKHX1_CV
XA9 CK_N CK_B AVDD AVSS AVDD AVSS IVX1_CV
XA10 DONE_N CK_A CK_N AVDD AVSS AVDD AVSS NDX1_CV
XA11 CK_SAMPLE DONE DONE_N AVDD AVSS AVDD AVSS NRX1_CV
XA12 CK_CMP CK_A AVDD AVSS AVDD AVSS IVX1_CV
XA13 AVDD AVSS TAPCELLB_CV
*XA14 DMY_CV
.ENDS


.SUBCKT SARMRYX1_CV CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 CMP_OP CMP_ON EN ENO RST_N AVDD AVSS AVDD AVSS SAREMX1_CV
XA2 ENO LCK_N AVDD AVSS AVDD AVSS IVX1_CV
XA4 CMP_OP CHL_OP RST_N EN LCK_N AVDD AVSS AVDD AVSS SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN LCK_N AVDD AVSS AVDD AVSS SARLTX1_CV
.ENDS

.SUBCKT SARDIGX1_CV CMP_OP CMP_ON EN RST_N ENO CP0 CP1 CN0 CN1 VREF AVDD AVSS
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS SARMRYX1_CV
XA2 CHL_ON CN1 VREF AVSS AVDD AVSS SWX2_CV
XA3 CN1 CP1 VREF AVSS AVDD AVSS SWX2_CV
XA4 CHL_OP CP0 VREF AVSS AVDD AVSS SWX2_CV
XA5 CP0 CN0 VREF AVSS AVDD AVSS SWX2_CV
XA6 AVDD AVSS TAPCELLB_CV
.ENDS

.SUBCKT SARDIGEX2_CV CMP_OP CMP_ON EN RST_N ENO DONE CP0 CP1 CN0 CN1 CEIN CEO CKS VREF AVDD AVSS
*XA0a DMY_CV
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON  AVDD AVSS SARMRYX1_CV

XA2 CHL_ON CN1 VREF AVSS AVDD AVSS SWX2_CV
XA3 CN1 CP1 VREF AVSS AVDD AVSS SWX2_CV
XA4 CHL_OP CP0 VREF AVSS AVDD AVSS SWX2_CV
XA5 CP0 CN0 VREF AVSS AVDD AVSS SWX2_CV

XA6 CN0 CP1 CE CKS AVDD AVSS AVDD AVSS SARCEX1_CV
XA7 ENO ENO_N AVDD AVSS AVDD AVSS IVX1_CV
XA8 ENO_N DONE AVDD AVSS AVDD AVSS IVX1_CV
XA9 ENO_N CE CE1 AVDD AVSS AVDD AVSS NDX1_CV
XA10 CE1 CE1_N AVDD AVSS AVDD AVSS IVX1_CV
XA11 CE1_N CEIN CEO1 AVDD AVSS AVDD AVSS NRX1_CV
XA12 CEO1 CEO AVDD AVSS AVDD AVSS IVX1_CV
XA13 AVDD AVSS TAPCELLB_CV
*XA14 DMY_CV
.ENDS

*-----------------------------------------------------------------------------
* SAR capacitors
*-----------------------------------------------------------------------------


.subckt CAP32C_CV C1A C1B C2 C4 C8 C16 CTOP AVSS
*XR1 CTOP NCa RM4
*XR2 AVSS Ncb RM4

XRES1A C1A NC1 RM1
XRES1B C1B NC2 RM1
XRES2 C2 NC3 RM1
XRES4 C4 NC4 RM1
XRES8 C8 NC5 RM1
XRES16 C16 NC6 RM1
.ends CAP32C_CV


*-----------------------------------------------------------------------------
* SAR CDACs
*-----------------------------------------------------------------------------


.SUBCKT CDAC7_CV   CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XC1  CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CTOP AVSS  CAP32C_CV
XC32a<0>  AVSS CP<0> CP<1> CP<2> CP<3> CP<7> CTOP AVSS  CAP32C_CV
X16ab       CP<5> CP<5> CP<5> CP<5> CP<4> CP<6> CTOP AVSS  CAP32C_CV
XC0  CP<9> CP<9> CP<9> CP<9> CP<9> CP<9> CTOP AVSS  CAP32C_CV
.ENDS CDAC7_CV

.SUBCKT CDAC8_CV  CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XC1  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CAP32C_CV
XC64a<0>  CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CTOP AVSS  CAP32C_CV
XC32a<0>  AVSS CP<0> CP<1> CP<2> CP<3> CP<7> CTOP AVSS  CAP32C_CV
XC128a<1>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CAP32C_CV 
XC128b<2>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CAP32C_CV
X16ab       CP<5> CP<5> CP<5> CP<5> CP<4> CP<6> CTOP AVSS  CAP32C_CV
XC64b<1>  CP<9> CP<9> CP<9> CP<9> CP<9> CP<9> CTOP AVSS  CAP32C_CV
XC0 CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CAP32C_CV
.ENDS CDAC8_CV

*-----------------------------------------------------------------------------
* SAR CDACs with logic
*-----------------------------------------------------------------------------

.SUBCKT SAR9B_CV_NOROUTE SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW  VREF AVDD AVSS

XB1  SAR_IP CK_SAMPLE_BSSW NCCA CEIN SARP SARN AVDD AVSS SARBSSW_CV
XB2  SAR_IN CK_SAMPLE_BSSW NCCB CEIN SARN SARP AVDD AVSS SARBSSW_CV


XDAC1  CP<11> CP<10>    D<7>  CP<8>  D<6>  CP<6>  D<5>  CP<4>  D<4>  D<3>  D<2>  D<1> SARP AVSS CDAC8_CV
XDAC2  D<8>   CN<10>    CN<9> CN<8>  CN<7> CN<6>  CN<5> CN<4>  CN<3> CN<2> CN<1> CN<0> SARN  AVSS CDAC8_CV

XA0 CMP_OP CMP_ON EN EN ENO0 DONE0   CP<10> CP<11> CN<10> D<8>  CEIN CEO0   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA1 CMP_OP CMP_ON ENO0 EN ENO1 DONE1 CP<8>  D<7>   CN<8>  CN<9> CEO0 CEO1   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA2 CMP_OP CMP_ON ENO1 EN ENO2 DONE2 CP<6>  D<6>   CN<6>  CN<7> CEO1 CEO2   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA3 CMP_OP CMP_ON ENO2 EN ENO3 DONE3 CP<4>  D<5>   CN<4>  CN<5> CEO2 CEO3   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA4 CMP_OP CMP_ON ENO3 EN ENO4 DONE4 NC2A   D<4>   CN<3>  NC2B  CEO3 CEO4   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA5 CMP_OP CMP_ON ENO4 EN ENO5 DONE5 NC3A   D<3>   CN<2>  NC3B  CEO4 CEO5   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA6 CMP_OP CMP_ON ENO5 EN ENO6 DONE6 NC4A   D<2>   CN<1>  NC4B  CEO5 CEO6   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA7 CMP_OP CMP_ON ENO6 EN ENO7 DONE7 NC5A   D<1>   CN<0>  NC5B  CEO6 CEO7   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA8 CMP_OP CMP_ON ENO7 EN ENO8 DONE  NC6A   D<0>   NC6C   NC6B  CEO7 CK_CMP CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV

XA20 SARP SARN CMP_OP CMP_ON CK_CMP CK_SAMPLE DONE AVDD AVSS SARCMPX1_CV
.ENDS


.SUBCKT SAR8B_CV SAR_IP SAR_IN SARN SARP DONE  D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW  VREF AVDD AVSS

XB1  SAR_IP CK_SAMPLE_BSSW NCCA CEIN SARP SARN AVDD AVSS SARBSSW_CV
XB2  SAR_IN CK_SAMPLE_BSSW NCCB CEIN SARN SARP AVDD AVSS SARBSSW_CV


XDAC1  CP<9>  CP<8>  D<6>  CP<6>  D<5>  CP<4>  D<4>  D<3>  D<2>  D<1> SARP AVSS CDAC7_CV
XDAC2  D<7> CN<8>  CN<7> CN<6>  CN<5> CN<4>  CN<3> CN<2> CN<1> CN<0> SARN  AVSS CDAC7_CV

*XA0 CMP_OP CMP_ON EN EN ENO0 DONE0   CP<10> CP<11> CN<10> D<8>  CEIN CEO0   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA0 CMP_OP CMP_ON EN EN ENO0 DONE0   CP<8>  CP<9>   CN<8>  D<7> CEIN CEO0   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA1 CMP_OP CMP_ON ENO0 EN ENO1 DONE1 CP<6>  D<6>   CN<6>  CN<7> CEO0 CEO1   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA2 CMP_OP CMP_ON ENO1 EN ENO2 DONE2 CP<4>  D<5>   CN<4>  CN<5> CEO1 CEO2   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA3 CMP_OP CMP_ON ENO2 EN ENO3 DONE3 NC2A   D<4>   CN<3>  NC2B  CEO2 CEO3   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA4 CMP_OP CMP_ON ENO3 EN ENO4 DONE4 NC3A   D<3>   CN<2>  NC3B  CEO3 CEO4   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA5 CMP_OP CMP_ON ENO4 EN ENO5 DONE5 NC4A   D<2>   CN<1>  NC4B  CEO4 CEO5   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA6 CMP_OP CMP_ON ENO5 EN ENO6 DONE6 NC5A   D<1>   CN<0>  NC5B  CEO5 CEO6   CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV
XA7 CMP_OP CMP_ON ENO6 EN ENO7 DONE  NC6A   D<0>   NC6C   NC6B  CEO6 CK_CMP CK_SAMPLE VREF AVDD AVSS SARDIGEX4_CV

XA20 SARP SARN CMP_OP CMP_ON CK_CMP CK_SAMPLE DONE AVDD AVSS SARCMPX1_CV
.ENDS

.subckt SARCAPTURE_CV CKS ENABLE CK_SAMPLE CK_SAMPLE_BSSW EN
+ D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0>
+ DO<7> DO<6> DO<5> DO<4> DO<3> DO<2> DO<1> DO<0>
+ DONE AVDD AVSS


XB07 D<7> DONE ENABLE_B DO<7> DN7 AVDD AVSS  DFRNQNX1_CV
XC08 D<6> DONE ENABLE_B DO<6> DN6 AVDD AVSS  DFRNQNX1_CV
XD09 D<5> DONE ENABLE_B DO<5> DN5 AVDD AVSS  DFRNQNX1_CV
XE10 D<4> DONE ENABLE_B DO<4> DN4 AVDD AVSS  DFRNQNX1_CV
XF11 D<3> DONE ENABLE_B DO<3> DN3 AVDD AVSS  DFRNQNX1_CV
XG12 D<2> DONE ENABLE_B DO<2> DN2 AVDD AVSS  DFRNQNX1_CV
XH13 D<1> DONE ENABLE_B DO<1> DN1 AVDD AVSS  DFRNQNX1_CV
XI14 D<0> DONE ENABLE_B DO<0> DM0 AVDD AVSS  DFRNQNX1_CV

XA1 AVDD AVSS TAPCELLB_CV
XA2 ENABLE ENABLE_N AVDD AVSS AVDD AVSS IVX1_CV
XA3 ENABLE_N ENABLE_B AVDD AVSS AVDD AVSS IVX1_CV
XA4 CKS CKS_B AVDD AVSS AVDD AVSS BFX1_CV
XA5 CKS_B ENABLE_N CK_SAMPLE AVDD AVSS AVDD AVSS ORX1_CV
XA5a CK_SAMPLE EN AVDD AVSS AVDD AVSS IVX1_CV
XA6 CKS_B ENABLE_B CK_SAMPLE_BSSW AVDD AVSS AVDD AVSS ANX1_CV
.ends


.subckt CAPT8B_CV CKS ENABLE CK_SAMPLE CK_SAMPLE_BSSW EN
+ D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0>
+ DO<7> DO<6> DO<5> DO<4> DO<3> DO<2> DO<1> DO<0>
+ DONE AVDD AVSS

XB07 D<7> DONE DO<7> DN7 AVDD AVSS  DFQNX1_CV
XC08 D<6> DONE DO<6> DN6 AVDD AVSS  DFQNX1_CV
XD09 D<5> DONE DO<5> DN5 AVDD AVSS  DFQNX1_CV
XE10 D<4> DONE DO<4> DN4 AVDD AVSS  DFQNX1_CV
XF11 D<3> DONE DO<3> DN3 AVDD AVSS  DFQNX1_CV
XG12 D<2> DONE DO<2> DN2 AVDD AVSS  DFQNX1_CV
XH13 D<1> DONE DO<1> DN1 AVDD AVSS  DFQNX1_CV
XI14 D<0> DONE DO<0> DM0 AVDD AVSS  DFQNX1_CV

XA1 AVDD AVSS TAPCELLB_CV
XA2 ENABLE ENABLE_N AVDD AVSS AVDD AVSS IVX1_CV
XA3 ENABLE_N ENABLE_B AVDD AVSS AVDD AVSS IVX1_CV
XA4 CKS CKS_B AVDD AVSS AVDD AVSS BFX1_CV
XA5 CKS_B ENABLE_N CK_SAMPLE AVDD AVSS AVDD AVSS ORX1_CV
XA5a CK_SAMPLE EN AVDD AVSS AVDD AVSS IVX1_CV
XA6 CKS_B ENABLE_B CK_SAMPLE_BSSW AVDD AVSS AVDD AVSS ANX1_CV
.ends
