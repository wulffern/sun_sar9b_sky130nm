magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 68 0 5702 13634
<< m1 >>
rect 1102 5166 1136 13600
rect 1102 5166 1136 13600
rect 1008 66 1042 13600
rect 1008 66 1042 13600
rect 914 10266 948 13600
rect 914 10266 948 13600
rect 820 1766 854 13600
rect 820 1766 854 13600
rect 726 3768 760 13600
rect 726 3768 760 13600
rect 632 8868 666 13600
rect 632 8868 666 13600
rect 538 8566 572 13600
rect 538 8566 572 13600
rect 444 9472 478 13600
rect 444 9472 478 13600
rect 350 4372 384 13600
rect 350 4372 384 13600
rect 256 4674 290 13600
rect 256 4674 290 13600
rect 162 4070 196 13600
rect 162 4070 196 13600
rect 68 4976 102 13600
rect 68 4976 102 13600
rect 1222 3466 1256 3558
rect 1222 3495 1378 3529
rect 1378 0 5668 34
<< m2 >>
rect 1136 5195 1222 5229
rect 1136 6705 1222 6739
rect 1136 5799 1222 5833
rect 1136 6403 1222 6437
rect 1136 6101 1222 6135
rect 1136 5497 1222 5531
rect 1136 11995 1222 12029
rect 1136 13505 1222 13539
rect 1136 12599 1222 12633
rect 1136 13203 1222 13237
rect 1136 12901 1222 12935
rect 1136 12297 1222 12331
rect 1042 95 1222 129
rect 1042 1605 1222 1639
rect 1042 699 1222 733
rect 1042 1303 1222 1337
rect 1042 1001 1222 1035
rect 1042 397 1222 431
rect 1042 6895 1222 6929
rect 1042 8405 1222 8439
rect 1042 7499 1222 7533
rect 1042 8103 1222 8137
rect 1042 7801 1222 7835
rect 1042 7197 1222 7231
rect 948 10295 1222 10329
rect 948 11805 1222 11839
rect 948 10899 1222 10933
rect 948 11503 1222 11537
rect 948 11201 1222 11235
rect 948 10597 1222 10631
rect 854 1795 1222 1829
rect 854 3305 1222 3339
rect 854 2399 1222 2433
rect 854 3003 1222 3037
rect 854 2701 1222 2735
rect 854 2097 1222 2131
rect 760 3797 1222 3831
rect 666 8897 1222 8931
rect 572 8595 1222 8629
rect 572 10105 1222 10139
rect 572 9199 1222 9233
rect 572 9803 1222 9837
rect 478 9501 1222 9535
rect 384 4401 1222 4435
rect 290 4703 1222 4737
rect 196 4099 1222 4133
rect 102 5005 1222 5039
<< locali >>
rect 1222 3466 1256 3558
<< viali >>
rect 1225 3472 1253 3500
rect 1225 3524 1253 3552
<< m3 >>
rect 1378 11900 1412 13634
use SUNSAR_CAP32C_CV XC1 
transform 1 0 1222 0 1 0
box 1222 0 5702 1700
use SUNSAR_CAP32C_CV XC64a<0> 
transform 1 0 1222 0 1 1700
box 1222 1700 5702 3400
use SUNSAR_CAP32C_CV XC32a<0> 
transform 1 0 1222 0 1 3400
box 1222 3400 5702 5100
use SUNSAR_CAP32C_CV XC128a<1> 
transform 1 0 1222 0 1 5100
box 1222 5100 5702 6800
use SUNSAR_CAP32C_CV XC128b<2> 
transform 1 0 1222 0 1 6800
box 1222 6800 5702 8500
use SUNSAR_CAP32C_CV X16ab 
transform 1 0 1222 0 1 8500
box 1222 8500 5702 10200
use SUNSAR_CAP32C_CV XC64b<1> 
transform 1 0 1222 0 1 10200
box 1222 10200 5702 11900
use SUNSAR_CAP32C_CV XC0 
transform 1 0 1222 0 1 11900
box 1222 11900 5702 13600
use SUNSAR_cut_M1M3_2x1 xcut0 
transform 1 0 1222 0 1 5195
box 1222 5195 1314 5229
use SUNSAR_cut_M2M3_1x2 xcut1 
transform 1 0 1102 0 1 5166
box 1102 5166 1136 5258
use SUNSAR_cut_M1M3_2x1 xcut2 
transform 1 0 1222 0 1 6705
box 1222 6705 1314 6739
use SUNSAR_cut_M2M3_1x2 xcut3 
transform 1 0 1102 0 1 6676
box 1102 6676 1136 6768
use SUNSAR_cut_M1M3_2x1 xcut4 
transform 1 0 1222 0 1 5799
box 1222 5799 1314 5833
use SUNSAR_cut_M2M3_1x2 xcut5 
transform 1 0 1102 0 1 5770
box 1102 5770 1136 5862
use SUNSAR_cut_M1M3_2x1 xcut6 
transform 1 0 1222 0 1 6403
box 1222 6403 1314 6437
use SUNSAR_cut_M2M3_1x2 xcut7 
transform 1 0 1102 0 1 6374
box 1102 6374 1136 6466
use SUNSAR_cut_M1M3_2x1 xcut8 
transform 1 0 1222 0 1 6101
box 1222 6101 1314 6135
use SUNSAR_cut_M2M3_1x2 xcut9 
transform 1 0 1102 0 1 6072
box 1102 6072 1136 6164
use SUNSAR_cut_M1M3_2x1 xcut10 
transform 1 0 1222 0 1 5497
box 1222 5497 1314 5531
use SUNSAR_cut_M2M3_1x2 xcut11 
transform 1 0 1102 0 1 5468
box 1102 5468 1136 5560
use SUNSAR_cut_M1M3_2x1 xcut12 
transform 1 0 1222 0 1 11995
box 1222 11995 1314 12029
use SUNSAR_cut_M2M3_1x2 xcut13 
transform 1 0 1102 0 1 11966
box 1102 11966 1136 12058
use SUNSAR_cut_M1M3_2x1 xcut14 
transform 1 0 1222 0 1 13505
box 1222 13505 1314 13539
use SUNSAR_cut_M2M3_1x2 xcut15 
transform 1 0 1102 0 1 13476
box 1102 13476 1136 13568
use SUNSAR_cut_M1M3_2x1 xcut16 
transform 1 0 1222 0 1 12599
box 1222 12599 1314 12633
use SUNSAR_cut_M2M3_1x2 xcut17 
transform 1 0 1102 0 1 12570
box 1102 12570 1136 12662
use SUNSAR_cut_M1M3_2x1 xcut18 
transform 1 0 1222 0 1 13203
box 1222 13203 1314 13237
use SUNSAR_cut_M2M3_1x2 xcut19 
transform 1 0 1102 0 1 13174
box 1102 13174 1136 13266
use SUNSAR_cut_M1M3_2x1 xcut20 
transform 1 0 1222 0 1 12901
box 1222 12901 1314 12935
use SUNSAR_cut_M2M3_1x2 xcut21 
transform 1 0 1102 0 1 12872
box 1102 12872 1136 12964
use SUNSAR_cut_M1M3_2x1 xcut22 
transform 1 0 1222 0 1 12297
box 1222 12297 1314 12331
use SUNSAR_cut_M2M3_1x2 xcut23 
transform 1 0 1102 0 1 12268
box 1102 12268 1136 12360
use SUNSAR_cut_M1M3_2x1 xcut24 
transform 1 0 1222 0 1 95
box 1222 95 1314 129
use SUNSAR_cut_M2M3_1x2 xcut25 
transform 1 0 1008 0 1 66
box 1008 66 1042 158
use SUNSAR_cut_M1M3_2x1 xcut26 
transform 1 0 1222 0 1 1605
box 1222 1605 1314 1639
use SUNSAR_cut_M2M3_1x2 xcut27 
transform 1 0 1008 0 1 1576
box 1008 1576 1042 1668
use SUNSAR_cut_M1M3_2x1 xcut28 
transform 1 0 1222 0 1 699
box 1222 699 1314 733
use SUNSAR_cut_M2M3_1x2 xcut29 
transform 1 0 1008 0 1 670
box 1008 670 1042 762
use SUNSAR_cut_M1M3_2x1 xcut30 
transform 1 0 1222 0 1 1303
box 1222 1303 1314 1337
use SUNSAR_cut_M2M3_1x2 xcut31 
transform 1 0 1008 0 1 1274
box 1008 1274 1042 1366
use SUNSAR_cut_M1M3_2x1 xcut32 
transform 1 0 1222 0 1 1001
box 1222 1001 1314 1035
use SUNSAR_cut_M2M3_1x2 xcut33 
transform 1 0 1008 0 1 972
box 1008 972 1042 1064
use SUNSAR_cut_M1M3_2x1 xcut34 
transform 1 0 1222 0 1 397
box 1222 397 1314 431
use SUNSAR_cut_M2M3_1x2 xcut35 
transform 1 0 1008 0 1 368
box 1008 368 1042 460
use SUNSAR_cut_M1M3_2x1 xcut36 
transform 1 0 1222 0 1 6895
box 1222 6895 1314 6929
use SUNSAR_cut_M2M3_1x2 xcut37 
transform 1 0 1008 0 1 6866
box 1008 6866 1042 6958
use SUNSAR_cut_M1M3_2x1 xcut38 
transform 1 0 1222 0 1 8405
box 1222 8405 1314 8439
use SUNSAR_cut_M2M3_1x2 xcut39 
transform 1 0 1008 0 1 8376
box 1008 8376 1042 8468
use SUNSAR_cut_M1M3_2x1 xcut40 
transform 1 0 1222 0 1 7499
box 1222 7499 1314 7533
use SUNSAR_cut_M2M3_1x2 xcut41 
transform 1 0 1008 0 1 7470
box 1008 7470 1042 7562
use SUNSAR_cut_M1M3_2x1 xcut42 
transform 1 0 1222 0 1 8103
box 1222 8103 1314 8137
use SUNSAR_cut_M2M3_1x2 xcut43 
transform 1 0 1008 0 1 8074
box 1008 8074 1042 8166
use SUNSAR_cut_M1M3_2x1 xcut44 
transform 1 0 1222 0 1 7801
box 1222 7801 1314 7835
use SUNSAR_cut_M2M3_1x2 xcut45 
transform 1 0 1008 0 1 7772
box 1008 7772 1042 7864
use SUNSAR_cut_M1M3_2x1 xcut46 
transform 1 0 1222 0 1 7197
box 1222 7197 1314 7231
use SUNSAR_cut_M2M3_1x2 xcut47 
transform 1 0 1008 0 1 7168
box 1008 7168 1042 7260
use SUNSAR_cut_M1M3_2x1 xcut48 
transform 1 0 1222 0 1 10295
box 1222 10295 1314 10329
use SUNSAR_cut_M2M3_1x2 xcut49 
transform 1 0 914 0 1 10266
box 914 10266 948 10358
use SUNSAR_cut_M1M3_2x1 xcut50 
transform 1 0 1222 0 1 11805
box 1222 11805 1314 11839
use SUNSAR_cut_M2M3_1x2 xcut51 
transform 1 0 914 0 1 11776
box 914 11776 948 11868
use SUNSAR_cut_M1M3_2x1 xcut52 
transform 1 0 1222 0 1 10899
box 1222 10899 1314 10933
use SUNSAR_cut_M2M3_1x2 xcut53 
transform 1 0 914 0 1 10870
box 914 10870 948 10962
use SUNSAR_cut_M1M3_2x1 xcut54 
transform 1 0 1222 0 1 11503
box 1222 11503 1314 11537
use SUNSAR_cut_M2M3_1x2 xcut55 
transform 1 0 914 0 1 11474
box 914 11474 948 11566
use SUNSAR_cut_M1M3_2x1 xcut56 
transform 1 0 1222 0 1 11201
box 1222 11201 1314 11235
use SUNSAR_cut_M2M3_1x2 xcut57 
transform 1 0 914 0 1 11172
box 914 11172 948 11264
use SUNSAR_cut_M1M3_2x1 xcut58 
transform 1 0 1222 0 1 10597
box 1222 10597 1314 10631
use SUNSAR_cut_M2M3_1x2 xcut59 
transform 1 0 914 0 1 10568
box 914 10568 948 10660
use SUNSAR_cut_M1M3_2x1 xcut60 
transform 1 0 1222 0 1 1795
box 1222 1795 1314 1829
use SUNSAR_cut_M2M3_1x2 xcut61 
transform 1 0 820 0 1 1766
box 820 1766 854 1858
use SUNSAR_cut_M1M3_2x1 xcut62 
transform 1 0 1222 0 1 3305
box 1222 3305 1314 3339
use SUNSAR_cut_M2M3_1x2 xcut63 
transform 1 0 820 0 1 3276
box 820 3276 854 3368
use SUNSAR_cut_M1M3_2x1 xcut64 
transform 1 0 1222 0 1 2399
box 1222 2399 1314 2433
use SUNSAR_cut_M2M3_1x2 xcut65 
transform 1 0 820 0 1 2370
box 820 2370 854 2462
use SUNSAR_cut_M1M3_2x1 xcut66 
transform 1 0 1222 0 1 3003
box 1222 3003 1314 3037
use SUNSAR_cut_M2M3_1x2 xcut67 
transform 1 0 820 0 1 2974
box 820 2974 854 3066
use SUNSAR_cut_M1M3_2x1 xcut68 
transform 1 0 1222 0 1 2701
box 1222 2701 1314 2735
use SUNSAR_cut_M2M3_1x2 xcut69 
transform 1 0 820 0 1 2672
box 820 2672 854 2764
use SUNSAR_cut_M1M3_2x1 xcut70 
transform 1 0 1222 0 1 2097
box 1222 2097 1314 2131
use SUNSAR_cut_M2M3_1x2 xcut71 
transform 1 0 820 0 1 2068
box 820 2068 854 2160
use SUNSAR_cut_M1M3_2x1 xcut72 
transform 1 0 1222 0 1 3797
box 1222 3797 1314 3831
use SUNSAR_cut_M2M3_1x2 xcut73 
transform 1 0 726 0 1 3768
box 726 3768 760 3860
use SUNSAR_cut_M1M3_2x1 xcut74 
transform 1 0 1222 0 1 8897
box 1222 8897 1314 8931
use SUNSAR_cut_M2M3_1x2 xcut75 
transform 1 0 632 0 1 8868
box 632 8868 666 8960
use SUNSAR_cut_M1M3_2x1 xcut76 
transform 1 0 1222 0 1 8595
box 1222 8595 1314 8629
use SUNSAR_cut_M2M3_1x2 xcut77 
transform 1 0 538 0 1 8566
box 538 8566 572 8658
use SUNSAR_cut_M1M3_2x1 xcut78 
transform 1 0 1222 0 1 10105
box 1222 10105 1314 10139
use SUNSAR_cut_M2M3_1x2 xcut79 
transform 1 0 538 0 1 10076
box 538 10076 572 10168
use SUNSAR_cut_M1M3_2x1 xcut80 
transform 1 0 1222 0 1 9199
box 1222 9199 1314 9233
use SUNSAR_cut_M2M3_1x2 xcut81 
transform 1 0 538 0 1 9170
box 538 9170 572 9262
use SUNSAR_cut_M1M3_2x1 xcut82 
transform 1 0 1222 0 1 9803
box 1222 9803 1314 9837
use SUNSAR_cut_M2M3_1x2 xcut83 
transform 1 0 538 0 1 9774
box 538 9774 572 9866
use SUNSAR_cut_M1M3_2x1 xcut84 
transform 1 0 1222 0 1 9501
box 1222 9501 1314 9535
use SUNSAR_cut_M2M3_1x2 xcut85 
transform 1 0 444 0 1 9472
box 444 9472 478 9564
use SUNSAR_cut_M1M3_2x1 xcut86 
transform 1 0 1222 0 1 4401
box 1222 4401 1314 4435
use SUNSAR_cut_M2M3_1x2 xcut87 
transform 1 0 350 0 1 4372
box 350 4372 384 4464
use SUNSAR_cut_M1M3_2x1 xcut88 
transform 1 0 1222 0 1 4703
box 1222 4703 1314 4737
use SUNSAR_cut_M2M3_1x2 xcut89 
transform 1 0 256 0 1 4674
box 256 4674 290 4766
use SUNSAR_cut_M1M3_2x1 xcut90 
transform 1 0 1222 0 1 4099
box 1222 4099 1314 4133
use SUNSAR_cut_M2M3_1x2 xcut91 
transform 1 0 162 0 1 4070
box 162 4070 196 4162
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 1222 0 1 5005
box 1222 5005 1314 5039
use SUNSAR_cut_M2M3_1x2 xcut93 
transform 1 0 68 0 1 4976
box 68 4976 102 5068
<< labels >>
flabel m1 s 1102 5166 1136 13600 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew signal bidirectional
flabel m1 s 1008 66 1042 13600 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew signal bidirectional
flabel m1 s 914 10266 948 13600 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew signal bidirectional
flabel m1 s 820 1766 854 13600 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew signal bidirectional
flabel m1 s 726 3768 760 13600 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew signal bidirectional
flabel m1 s 632 8868 666 13600 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew signal bidirectional
flabel m1 s 538 8566 572 13600 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew signal bidirectional
flabel m1 s 444 9472 478 13600 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew signal bidirectional
flabel m1 s 350 4372 384 13600 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew signal bidirectional
flabel m1 s 256 4674 290 13600 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew signal bidirectional
flabel m1 s 162 4070 196 13600 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew signal bidirectional
flabel m1 s 68 4976 102 13600 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew signal bidirectional
flabel m1 s 1378 0 5668 34 0 FreeSans 400 0 0 0 AVSS
port 14 nsew signal bidirectional
flabel m3 s 1378 11900 1412 13634 0 FreeSans 400 0 0 0 CTOP
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 68 0 5702 13634
<< end >>
