magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect -961 -932 12139 18531
<< m3 >>
rect 4290 9572 11220 9606
rect 4290 9758 11220 9792
rect 10161 9928 10195 12770
rect 10299 9928 10333 15058
rect 97 9978 131 14354
rect 97 9978 131 14354
rect 2169 10071 2203 14354
rect 2617 10164 2651 14354
rect 442 10257 476 14369
rect 1881 10350 1915 14369
rect 1881 10350 1915 14369
rect 2962 10443 2996 14369
rect 2962 10443 2996 14369
rect 4401 10536 4435 14369
rect 4401 10536 4435 14369
rect 5482 10629 5516 14369
rect 5482 10629 5516 14369
rect 6921 10722 6955 14369
rect 6921 10722 6955 14369
rect 8002 10815 8036 14369
rect 8002 10815 8036 14369
rect 513 10908 547 14809
rect 1810 11001 1844 14809
rect 3033 11094 3067 14809
rect 592 11187 626 15249
rect 1732 11280 1766 15249
rect 3112 11373 3146 15249
rect 4252 11466 4286 15249
rect 5632 11559 5666 15249
rect 6772 11652 6806 15249
rect 8152 11745 8186 15249
rect 297 12083 389 17811
rect 1969 12083 2061 17811
rect 2817 12083 2909 17811
rect 4489 12083 4581 17811
rect 5337 12083 5429 17811
rect 7009 12083 7101 17811
rect 7857 12083 7949 17811
rect 9529 12083 9621 17811
rect 10377 12083 10469 17811
rect 4399 -360 4491 2400
rect 6687 -360 6779 2400
rect 693 12083 785 18171
rect 1573 12083 1665 18171
rect 3213 12083 3305 18171
rect 4093 12083 4185 18171
rect 5733 12083 5825 18171
rect 6613 12083 6705 18171
rect 8253 12083 8345 18171
rect 9133 12083 9225 18171
rect 10773 12083 10865 18171
rect 4003 -720 4095 2400
rect 7083 -720 7175 2400
rect 981 14046 1073 18531
rect 1285 14046 1377 18531
rect 3501 14046 3593 18531
rect 3805 14046 3897 18531
rect 6021 14046 6113 18531
rect 6325 14046 6417 18531
rect 8541 14046 8633 18531
rect 8845 14046 8937 18531
rect 4688 -932 4722 1469
rect 6456 -932 6490 1469
rect 4937 555 5157 589
rect 4307 2493 4937 2527
rect 6021 555 6207 589
rect 6207 2493 6871 2527
rect 5157 555 5241 589
rect 5241 1259 6021 1293
rect 5241 555 5275 1293
rect 5103 115 5195 149
rect 5983 115 6075 149
rect 9441 14369 9475 14461
<< m2 >>
rect 6854 9327 6888 9606
rect 4290 9327 4324 9792
rect 97 9944 6612 9978
rect 2169 10037 6424 10071
rect 2617 10130 6236 10164
rect 442 10223 4600 10257
rect 1881 10316 4788 10350
rect 2962 10409 4976 10443
rect 4401 10502 5164 10536
rect 5224 10595 5516 10629
rect 5318 10688 6955 10722
rect 5412 10781 8036 10815
rect 513 10874 4694 10908
rect 1810 10967 4882 11001
rect 3033 11060 5070 11094
rect 592 11153 6518 11187
rect 1732 11246 6330 11280
rect 3112 11339 6142 11373
rect 4252 11432 6048 11466
rect 5632 11525 5954 11559
rect 5826 11618 6806 11652
rect 5732 11711 8186 11745
rect 4636 -826 4670 281
rect 6508 -826 6542 281
rect -927 16994 81 17028
rect 693 17231 861 17265
rect 861 16930 2169 16964
rect 2135 16930 2169 17028
rect 861 16930 895 17265
rect 3213 17231 3381 17265
rect 3381 16930 4689 16964
rect 4655 16930 4689 17028
rect 3381 16930 3415 17265
rect 5733 17231 5901 17265
rect 5901 16930 7209 16964
rect 7175 16930 7209 17028
rect 5901 16930 5935 17265
rect 8253 17231 8421 17265
rect 8421 16930 9729 16964
rect 9695 16930 9729 17028
rect 8421 16930 8455 17265
rect 81 15698 9837 15732
rect 47 15698 81 15796
rect 2135 15698 2169 15796
rect 2567 15698 2601 15796
rect 4655 15698 4689 15796
rect 5087 15698 5121 15796
rect 7175 15698 7209 15796
rect 7607 15698 7641 15796
rect 9695 15698 9729 15796
rect 709 12462 861 12496
rect 861 12266 2169 12300
rect 2135 12266 2169 12364
rect 861 12266 895 12496
rect 3229 12462 3381 12496
rect 3381 12266 4689 12300
rect 4655 12266 4689 12364
rect 3381 12266 3415 12496
rect 5749 12462 5901 12496
rect 5901 12266 7209 12300
rect 7175 12266 7209 12364
rect 5901 12266 5935 12496
rect 8269 12462 8421 12496
rect 8421 12266 9729 12300
rect 9695 12266 9729 12364
rect 8421 12266 8455 12496
rect 1557 12462 1709 12496
rect 1709 12462 1743 12526
rect 1709 12526 2617 12560
rect 2583 12330 2617 12560
rect 4077 12462 4229 12496
rect 4229 12462 4263 12526
rect 4229 12526 5137 12560
rect 5103 12330 5137 12560
rect 6597 12462 6749 12496
rect 6749 12462 6783 12526
rect 6749 12526 7657 12560
rect 7623 12330 7657 12560
rect 9117 12462 9269 12496
rect 9269 12462 9303 12526
rect 97 13348 9821 13382
rect 63 13210 97 13382
rect 2135 13210 2169 13382
rect 2583 13210 2617 13382
rect 4655 13210 4689 13382
rect 5103 13210 5137 13382
rect 7175 13210 7209 13382
rect 7623 13210 7657 13382
rect 9695 13210 9729 13382
rect 81 13424 9837 13458
rect 47 13424 81 13596
rect 2135 13424 2169 13596
rect 2567 13424 2601 13596
rect 4655 13424 4689 13596
rect 5087 13424 5121 13596
rect 7175 13424 7209 13596
rect 7607 13424 7641 13596
rect 9695 13424 9729 13596
rect 189 13738 909 13772
rect 909 13738 1449 13772
rect 909 13738 3537 13772
rect 909 13738 3969 13772
rect 909 13738 6057 13772
rect 909 13738 6489 13772
rect 909 13738 8577 13772
rect 909 13738 9009 13772
rect 351 16334 435 16368
rect 435 16334 469 16368
rect 2007 16334 2091 16368
rect 2091 16334 2125 16368
rect 2871 16334 2955 16368
rect 2955 16334 2989 16368
rect 4527 16334 4611 16368
rect 4611 16334 4645 16368
rect 5391 16334 5475 16368
rect 5475 16334 5509 16368
rect 7047 16334 7131 16368
rect 7131 16334 7165 16368
rect 7911 16334 7995 16368
rect 7995 16334 8029 16368
rect 9567 16334 9651 16368
rect 9651 16554 10215 16588
rect 9651 16334 9685 16588
rect 10103 13799 10431 13833
rect 9791 13244 10103 13278
rect 10103 13244 10137 13833
rect 9775 13210 9821 13244
rect 9783 13562 9867 13596
rect 9867 14256 10803 14290
rect 9867 13562 9901 14290
rect 10773 14222 10827 14256
rect 11043 16466 11127 16500
rect 9807 15904 11127 15938
rect 11127 15904 11161 16500
rect 9783 15938 9837 15972
rect 9171 17214 9933 17248
rect 9933 16747 10215 16781
rect 9933 16747 9967 17248
rect 5157 1259 5241 1293
rect 5241 555 6021 589
rect 5241 555 5275 1293
rect 81 13738 1017 13772
<< m4 >>
rect 10161 9758 10195 9928
rect 10299 9572 10333 9928
rect 4937 555 4971 2527
rect 6207 555 6241 2527
<< m1 >>
rect 6578 9293 6612 9944
rect 6390 9293 6424 10037
rect 6202 9293 6236 10130
rect 4566 9293 4600 10223
rect 4754 9293 4788 10316
rect 4942 9293 4976 10409
rect 5130 9293 5164 10502
rect 5224 9293 5258 10595
rect 5318 9293 5352 10688
rect 5412 9293 5446 10781
rect 4660 9293 4694 10874
rect 4848 9293 4882 10967
rect 5036 9293 5070 11060
rect 6484 9293 6518 11153
rect 6296 9293 6330 11246
rect 6108 9293 6142 11339
rect 6014 9293 6048 11432
rect 5920 9293 5954 11525
rect 5826 9293 5860 11618
rect 5732 9293 5766 11711
rect 11581 -360 11673 17811
rect -495 -360 11673 -268
rect -495 17719 11673 17811
rect -495 -360 -403 17811
rect 11581 -360 11673 17811
rect 11941 -720 12033 18171
rect -855 -720 12033 -628
rect -855 18079 12033 18171
rect -855 -720 -763 18171
rect 11941 -720 12033 18171
rect -855 18439 12033 18531
rect -855 18439 12033 18531
rect 12105 -826 12139 18531
rect -855 -826 12139 -792
rect 12105 -826 12139 18531
rect -961 -932 12139 -898
rect -961 -932 -927 18531
rect 1557 17214 1725 17248
rect 1725 16930 2601 16964
rect 2567 16930 2601 17028
rect 1725 16930 1759 17248
rect 4077 17214 4245 17248
rect 4245 16930 5121 16964
rect 5087 16930 5121 17028
rect 4245 16930 4279 17248
rect 6597 17214 6765 17248
rect 6765 16930 7641 16964
rect 7607 16930 7641 17028
rect 6765 16930 6799 17248
rect -495 2493 34 2527
rect -495 4193 34 4227
rect -495 5893 34 5927
rect -495 7593 34 7627
rect 11144 2493 11673 2527
rect 11144 4193 11673 4227
rect 11144 5893 11673 5927
rect 11144 7593 11673 7627
<< locali >>
rect 9513 16334 9621 16368
rect 81 15762 189 15796
rect 909 13738 1017 13772
rect 5103 1259 5211 1293
rect 5103 555 5211 589
use SUNSAR_SARBSSW_CV XB1 
transform -1 0 5589 0 1 0
box 5589 0 11313 2400
use SUNSAR_SARBSSW_CV XB2 
transform 1 0 5589 0 1 0
box 5589 0 11313 2400
use SUNSAR_CDAC7_CV XDAC1 
transform -1 0 5514 0 1 2493
box 5514 2493 10960 9327
use SUNSAR_CDAC7_CV XDAC2 
transform 1 0 5664 0 1 2493
box 5664 2493 11110 9327
use SUNSAR_SARDIGEX4_CV XA0 
transform 1 0 -81 0 1 12083
box -81 12083 1179 17451
use SUNSAR_SARDIGEX4_CV XA1 
transform -1 0 2439 0 1 12083
box 2439 12083 3699 17451
use SUNSAR_SARDIGEX4_CV XA2 
transform 1 0 2439 0 1 12083
box 2439 12083 3699 17451
use SUNSAR_SARDIGEX4_CV XA3 
transform -1 0 4959 0 1 12083
box 4959 12083 6219 17451
use SUNSAR_SARDIGEX4_CV XA4 
transform 1 0 4959 0 1 12083
box 4959 12083 6219 17451
use SUNSAR_SARDIGEX4_CV XA5 
transform -1 0 7479 0 1 12083
box 7479 12083 8739 17451
use SUNSAR_SARDIGEX4_CV XA6 
transform 1 0 7479 0 1 12083
box 7479 12083 8739 17451
use SUNSAR_SARDIGEX4_CV XA7 
transform -1 0 9999 0 1 12083
box 9999 12083 11259 17451
use SUNSAR_SARCMPX1_CV XA20 
transform 1 0 9999 0 1 12083
box 9999 12083 11259 17011
use SUNSAR_cut_M3M4_1x2 xcut0 
transform 1 0 6854 0 1 9327
box 6854 9327 6888 9419
use SUNSAR_cut_M3M4_2x1 xcut1 
transform 1 0 6854 0 1 9572
box 6854 9572 6946 9606
use SUNSAR_cut_M3M4_1x2 xcut2 
transform 1 0 4290 0 1 9327
box 4290 9327 4324 9419
use SUNSAR_cut_M3M4_2x1 xcut3 
transform 1 0 4290 0 1 9758
box 4290 9758 4382 9792
use SUNSAR_cut_M2M4_2x1 xcut4 
transform 1 0 10161 0 1 12770
box 10161 12770 10253 12804
use SUNSAR_cut_M4M5_2x1 xcut5 
transform 1 0 10161 0 1 9758
box 10161 9758 10257 9792
use SUNSAR_cut_M4M5_1x2 xcut6 
transform 1 0 10161 0 1 9928
box 10161 9928 10195 10024
use SUNSAR_cut_M3M4_2x1 xcut7 
transform 1 0 10241 0 1 15058
box 10241 15058 10333 15092
use SUNSAR_cut_M2M3_2x1 xcut8 
transform 1 0 10161 0 1 15058
box 10161 15058 10253 15092
use SUNSAR_cut_M4M5_2x1 xcut9 
transform 1 0 10299 0 1 9572
box 10299 9572 10395 9606
use SUNSAR_cut_M4M5_1x2 xcut10 
transform 1 0 10299 0 1 9928
box 10299 9928 10333 10024
use SUNSAR_cut_M3M4_1x2 xcut11 
transform 1 0 97 0 1 9915
box 97 9915 131 10007
use SUNSAR_cut_M2M3_1x2 xcut12 
transform 1 0 6578 0 1 9915
box 6578 9915 6612 10007
use SUNSAR_cut_M3M4_1x2 xcut13 
transform 1 0 2169 0 1 10008
box 2169 10008 2203 10100
use SUNSAR_cut_M2M3_1x2 xcut14 
transform 1 0 6390 0 1 10008
box 6390 10008 6424 10100
use SUNSAR_cut_M3M4_1x2 xcut15 
transform 1 0 2617 0 1 10101
box 2617 10101 2651 10193
use SUNSAR_cut_M2M3_1x2 xcut16 
transform 1 0 6202 0 1 10101
box 6202 10101 6236 10193
use SUNSAR_cut_M3M4_1x2 xcut17 
transform 1 0 442 0 1 10194
box 442 10194 476 10286
use SUNSAR_cut_M2M3_1x2 xcut18 
transform 1 0 4566 0 1 10194
box 4566 10194 4600 10286
use SUNSAR_cut_M3M4_1x2 xcut19 
transform 1 0 1881 0 1 10287
box 1881 10287 1915 10379
use SUNSAR_cut_M2M3_1x2 xcut20 
transform 1 0 4754 0 1 10287
box 4754 10287 4788 10379
use SUNSAR_cut_M3M4_1x2 xcut21 
transform 1 0 2962 0 1 10380
box 2962 10380 2996 10472
use SUNSAR_cut_M2M3_1x2 xcut22 
transform 1 0 4942 0 1 10380
box 4942 10380 4976 10472
use SUNSAR_cut_M3M4_1x2 xcut23 
transform 1 0 4401 0 1 10473
box 4401 10473 4435 10565
use SUNSAR_cut_M2M3_1x2 xcut24 
transform 1 0 5130 0 1 10473
box 5130 10473 5164 10565
use SUNSAR_cut_M3M4_1x2 xcut25 
transform 1 0 5482 0 1 10566
box 5482 10566 5516 10658
use SUNSAR_cut_M2M3_1x2 xcut26 
transform 1 0 5224 0 1 10566
box 5224 10566 5258 10658
use SUNSAR_cut_M3M4_1x2 xcut27 
transform 1 0 6921 0 1 10659
box 6921 10659 6955 10751
use SUNSAR_cut_M2M3_1x2 xcut28 
transform 1 0 5318 0 1 10659
box 5318 10659 5352 10751
use SUNSAR_cut_M3M4_1x2 xcut29 
transform 1 0 8002 0 1 10752
box 8002 10752 8036 10844
use SUNSAR_cut_M2M3_1x2 xcut30 
transform 1 0 5412 0 1 10752
box 5412 10752 5446 10844
use SUNSAR_cut_M3M4_1x2 xcut31 
transform 1 0 513 0 1 10845
box 513 10845 547 10937
use SUNSAR_cut_M2M3_1x2 xcut32 
transform 1 0 4660 0 1 10845
box 4660 10845 4694 10937
use SUNSAR_cut_M3M4_1x2 xcut33 
transform 1 0 1810 0 1 10938
box 1810 10938 1844 11030
use SUNSAR_cut_M2M3_1x2 xcut34 
transform 1 0 4848 0 1 10938
box 4848 10938 4882 11030
use SUNSAR_cut_M3M4_1x2 xcut35 
transform 1 0 3033 0 1 11031
box 3033 11031 3067 11123
use SUNSAR_cut_M2M3_1x2 xcut36 
transform 1 0 5036 0 1 11031
box 5036 11031 5070 11123
use SUNSAR_cut_M3M4_1x2 xcut37 
transform 1 0 592 0 1 11124
box 592 11124 626 11216
use SUNSAR_cut_M2M3_1x2 xcut38 
transform 1 0 6484 0 1 11124
box 6484 11124 6518 11216
use SUNSAR_cut_M3M4_1x2 xcut39 
transform 1 0 1732 0 1 11217
box 1732 11217 1766 11309
use SUNSAR_cut_M2M3_1x2 xcut40 
transform 1 0 6296 0 1 11217
box 6296 11217 6330 11309
use SUNSAR_cut_M3M4_1x2 xcut41 
transform 1 0 3112 0 1 11310
box 3112 11310 3146 11402
use SUNSAR_cut_M2M3_1x2 xcut42 
transform 1 0 6108 0 1 11310
box 6108 11310 6142 11402
use SUNSAR_cut_M3M4_1x2 xcut43 
transform 1 0 4252 0 1 11403
box 4252 11403 4286 11495
use SUNSAR_cut_M2M3_1x2 xcut44 
transform 1 0 6014 0 1 11403
box 6014 11403 6048 11495
use SUNSAR_cut_M3M4_1x2 xcut45 
transform 1 0 5632 0 1 11496
box 5632 11496 5666 11588
use SUNSAR_cut_M2M3_1x2 xcut46 
transform 1 0 5920 0 1 11496
box 5920 11496 5954 11588
use SUNSAR_cut_M3M4_1x2 xcut47 
transform 1 0 6772 0 1 11589
box 6772 11589 6806 11681
use SUNSAR_cut_M2M3_1x2 xcut48 
transform 1 0 5826 0 1 11589
box 5826 11589 5860 11681
use SUNSAR_cut_M3M4_1x2 xcut49 
transform 1 0 8152 0 1 11682
box 8152 11682 8186 11774
use SUNSAR_cut_M2M3_1x2 xcut50 
transform 1 0 5732 0 1 11682
box 5732 11682 5766 11774
use SUNSAR_cut_M2M4_2x2 xcut51 
transform 1 0 297 0 1 17719
box 297 17719 389 17811
use SUNSAR_cut_M2M4_2x2 xcut52 
transform 1 0 1969 0 1 17719
box 1969 17719 2061 17811
use SUNSAR_cut_M2M4_2x2 xcut53 
transform 1 0 2817 0 1 17719
box 2817 17719 2909 17811
use SUNSAR_cut_M2M4_2x2 xcut54 
transform 1 0 4489 0 1 17719
box 4489 17719 4581 17811
use SUNSAR_cut_M2M4_2x2 xcut55 
transform 1 0 5337 0 1 17719
box 5337 17719 5429 17811
use SUNSAR_cut_M2M4_2x2 xcut56 
transform 1 0 7009 0 1 17719
box 7009 17719 7101 17811
use SUNSAR_cut_M2M4_2x2 xcut57 
transform 1 0 7857 0 1 17719
box 7857 17719 7949 17811
use SUNSAR_cut_M2M4_2x2 xcut58 
transform 1 0 9529 0 1 17719
box 9529 17719 9621 17811
use SUNSAR_cut_M2M4_2x2 xcut59 
transform 1 0 10377 0 1 17719
box 10377 17719 10469 17811
use SUNSAR_cut_M2M4_2x2 xcut60 
transform 1 0 4399 0 1 -360
box 4399 -360 4491 -268
use SUNSAR_cut_M2M4_2x2 xcut61 
transform 1 0 6687 0 1 -360
box 6687 -360 6779 -268
use SUNSAR_cut_M2M4_2x2 xcut62 
transform 1 0 693 0 1 18079
box 693 18079 785 18171
use SUNSAR_cut_M2M4_2x2 xcut63 
transform 1 0 1573 0 1 18079
box 1573 18079 1665 18171
use SUNSAR_cut_M2M4_2x2 xcut64 
transform 1 0 3213 0 1 18079
box 3213 18079 3305 18171
use SUNSAR_cut_M2M4_2x2 xcut65 
transform 1 0 4093 0 1 18079
box 4093 18079 4185 18171
use SUNSAR_cut_M2M4_2x2 xcut66 
transform 1 0 5733 0 1 18079
box 5733 18079 5825 18171
use SUNSAR_cut_M2M4_2x2 xcut67 
transform 1 0 6613 0 1 18079
box 6613 18079 6705 18171
use SUNSAR_cut_M2M4_2x2 xcut68 
transform 1 0 8253 0 1 18079
box 8253 18079 8345 18171
use SUNSAR_cut_M2M4_2x2 xcut69 
transform 1 0 9133 0 1 18079
box 9133 18079 9225 18171
use SUNSAR_cut_M2M4_2x2 xcut70 
transform 1 0 10773 0 1 18079
box 10773 18079 10865 18171
use SUNSAR_cut_M2M4_2x2 xcut71 
transform 1 0 4003 0 1 -720
box 4003 -720 4095 -628
use SUNSAR_cut_M2M4_2x2 xcut72 
transform 1 0 7083 0 1 -720
box 7083 -720 7175 -628
use SUNSAR_cut_M2M4_2x2 xcut73 
transform 1 0 981 0 1 18439
box 981 18439 1073 18531
use SUNSAR_cut_M2M4_2x2 xcut74 
transform 1 0 1285 0 1 18439
box 1285 18439 1377 18531
use SUNSAR_cut_M2M4_2x2 xcut75 
transform 1 0 3501 0 1 18439
box 3501 18439 3593 18531
use SUNSAR_cut_M2M4_2x2 xcut76 
transform 1 0 3805 0 1 18439
box 3805 18439 3897 18531
use SUNSAR_cut_M2M4_2x2 xcut77 
transform 1 0 6021 0 1 18439
box 6021 18439 6113 18531
use SUNSAR_cut_M2M4_2x2 xcut78 
transform 1 0 6325 0 1 18439
box 6325 18439 6417 18531
use SUNSAR_cut_M2M4_2x2 xcut79 
transform 1 0 8541 0 1 18439
box 8541 18439 8633 18531
use SUNSAR_cut_M2M4_2x2 xcut80 
transform 1 0 8845 0 1 18439
box 8845 18439 8937 18531
use SUNSAR_cut_M1M3_2x1 xcut81 
transform 1 0 4607 0 1 247
box 4607 247 4699 281
use SUNSAR_cut_M2M3_2x1 xcut82 
transform 1 0 4607 0 1 -826
box 4607 -826 4699 -792
use SUNSAR_cut_M1M3_2x1 xcut83 
transform 1 0 6479 0 1 247
box 6479 247 6571 281
use SUNSAR_cut_M2M3_2x1 xcut84 
transform 1 0 6479 0 1 -826
box 6479 -826 6571 -792
use SUNSAR_cut_M1M3_2x1 xcut85 
transform 1 0 81 0 1 16994
box 81 16994 173 17028
use SUNSAR_cut_M2M3_1x2 xcut86 
transform 1 0 -961 0 1 16965
box -961 16965 -927 17057
use SUNSAR_cut_M2M4_2x1 xcut87 
transform 1 0 4659 0 1 -932
box 4659 -932 4751 -898
use SUNSAR_cut_M2M4_2x1 xcut88 
transform 1 0 6427 0 1 -932
box 6427 -932 6519 -898
use SUNSAR_cut_M1M3_2x1 xcut89 
transform 1 0 693 0 1 17231
box 693 17231 785 17265
use SUNSAR_cut_M1M3_2x1 xcut90 
transform 1 0 2169 0 1 16994
box 2169 16994 2261 17028
use SUNSAR_cut_M1M3_2x1 xcut91 
transform 1 0 3213 0 1 17231
box 3213 17231 3305 17265
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 4689 0 1 16994
box 4689 16994 4781 17028
use SUNSAR_cut_M1M3_2x1 xcut93 
transform 1 0 5733 0 1 17231
box 5733 17231 5825 17265
use SUNSAR_cut_M1M3_2x1 xcut94 
transform 1 0 7209 0 1 16994
box 7209 16994 7301 17028
use SUNSAR_cut_M1M3_2x1 xcut95 
transform 1 0 8253 0 1 17231
box 8253 17231 8345 17265
use SUNSAR_cut_M1M3_2x1 xcut96 
transform 1 0 9729 0 1 16994
box 9729 16994 9821 17028
use SUNSAR_cut_M1M3_2x1 xcut97 
transform 1 0 81 0 1 15762
box 81 15762 173 15796
use SUNSAR_cut_M1M3_2x1 xcut98 
transform 1 0 2169 0 1 15762
box 2169 15762 2261 15796
use SUNSAR_cut_M1M3_2x1 xcut99 
transform 1 0 2601 0 1 15762
box 2601 15762 2693 15796
use SUNSAR_cut_M1M3_2x1 xcut100 
transform 1 0 4689 0 1 15762
box 4689 15762 4781 15796
use SUNSAR_cut_M1M3_2x1 xcut101 
transform 1 0 5121 0 1 15762
box 5121 15762 5213 15796
use SUNSAR_cut_M1M3_2x1 xcut102 
transform 1 0 7209 0 1 15762
box 7209 15762 7301 15796
use SUNSAR_cut_M1M3_2x1 xcut103 
transform 1 0 7641 0 1 15762
box 7641 15762 7733 15796
use SUNSAR_cut_M1M3_2x1 xcut104 
transform 1 0 9729 0 1 15762
box 9729 15762 9821 15796
use SUNSAR_cut_M1M2_2x1 xcut105 
transform 1 0 1557 0 1 17214
box 1557 17214 1649 17248
use SUNSAR_cut_M1M2_2x1 xcut106 
transform 1 0 2601 0 1 16994
box 2601 16994 2693 17028
use SUNSAR_cut_M1M2_2x1 xcut107 
transform 1 0 4077 0 1 17214
box 4077 17214 4169 17248
use SUNSAR_cut_M1M2_2x1 xcut108 
transform 1 0 5121 0 1 16994
box 5121 16994 5213 17028
use SUNSAR_cut_M1M2_2x1 xcut109 
transform 1 0 6597 0 1 17214
box 6597 17214 6689 17248
use SUNSAR_cut_M1M2_2x1 xcut110 
transform 1 0 7641 0 1 16994
box 7641 16994 7733 17028
use SUNSAR_cut_M1M3_2x1 xcut111 
transform 1 0 81 0 1 13562
box 81 13562 173 13596
use SUNSAR_cut_M1M3_2x1 xcut112 
transform 1 0 2169 0 1 13562
box 2169 13562 2261 13596
use SUNSAR_cut_M1M3_2x1 xcut113 
transform 1 0 2601 0 1 13562
box 2601 13562 2693 13596
use SUNSAR_cut_M1M3_2x1 xcut114 
transform 1 0 4689 0 1 13562
box 4689 13562 4781 13596
use SUNSAR_cut_M1M3_2x1 xcut115 
transform 1 0 5121 0 1 13562
box 5121 13562 5213 13596
use SUNSAR_cut_M1M3_2x1 xcut116 
transform 1 0 7209 0 1 13562
box 7209 13562 7301 13596
use SUNSAR_cut_M1M3_2x1 xcut117 
transform 1 0 7641 0 1 13562
box 7641 13562 7733 13596
use SUNSAR_cut_M1M3_2x1 xcut118 
transform 1 0 9729 0 1 13562
box 9729 13562 9821 13596
use SUNSAR_cut_M1M3_2x1 xcut119 
transform 1 0 909 0 1 13738
box 909 13738 1001 13772
use SUNSAR_cut_M1M3_2x1 xcut120 
transform 1 0 1341 0 1 13738
box 1341 13738 1433 13772
use SUNSAR_cut_M1M3_2x1 xcut121 
transform 1 0 3429 0 1 13738
box 3429 13738 3521 13772
use SUNSAR_cut_M1M3_2x1 xcut122 
transform 1 0 3861 0 1 13738
box 3861 13738 3953 13772
use SUNSAR_cut_M1M3_2x1 xcut123 
transform 1 0 5949 0 1 13738
box 5949 13738 6041 13772
use SUNSAR_cut_M1M3_2x1 xcut124 
transform 1 0 6381 0 1 13738
box 6381 13738 6473 13772
use SUNSAR_cut_M1M3_2x1 xcut125 
transform 1 0 8469 0 1 13738
box 8469 13738 8561 13772
use SUNSAR_cut_M1M3_2x1 xcut126 
transform 1 0 8901 0 1 13738
box 8901 13738 8993 13772
use SUNSAR_cut_M1M3_2x1 xcut127 
transform 1 0 297 0 1 16334
box 297 16334 389 16368
use SUNSAR_cut_M1M3_2x1 xcut128 
transform 1 0 1953 0 1 16334
box 1953 16334 2045 16368
use SUNSAR_cut_M1M3_2x1 xcut129 
transform 1 0 2817 0 1 16334
box 2817 16334 2909 16368
use SUNSAR_cut_M1M3_2x1 xcut130 
transform 1 0 4473 0 1 16334
box 4473 16334 4565 16368
use SUNSAR_cut_M1M3_2x1 xcut131 
transform 1 0 5337 0 1 16334
box 5337 16334 5429 16368
use SUNSAR_cut_M1M3_2x1 xcut132 
transform 1 0 6993 0 1 16334
box 6993 16334 7085 16368
use SUNSAR_cut_M1M3_2x1 xcut133 
transform 1 0 7857 0 1 16334
box 7857 16334 7949 16368
use SUNSAR_cut_M1M3_2x1 xcut134 
transform 1 0 9513 0 1 16334
box 9513 16334 9605 16368
use SUNSAR_cut_M1M3_2x1 xcut135 
transform 1 0 10161 0 1 16554
box 10161 16554 10253 16588
use SUNSAR_cut_M1M3_2x1 xcut136 
transform 1 0 10393 0 1 13799
box 10393 13799 10485 13833
use SUNSAR_cut_M1M3_2x1 xcut137 
transform 1 0 10773 0 1 14222
box 10773 14222 10865 14256
use SUNSAR_cut_M1M3_2x1 xcut138 
transform 1 0 10989 0 1 16466
box 10989 16466 11081 16500
use SUNSAR_cut_M1M3_2x1 xcut139 
transform 1 0 9729 0 1 15938
box 9729 15938 9821 15972
use SUNSAR_cut_M1M3_2x1 xcut140 
transform 1 0 9117 0 1 17214
box 9117 17214 9209 17248
use SUNSAR_cut_M1M3_2x1 xcut141 
transform 1 0 10161 0 1 16747
box 10161 16747 10253 16781
use SUNSAR_cut_M4M5_1x2 xcut142 
transform 1 0 4937 0 1 555
box 4937 555 4971 651
use SUNSAR_cut_M4M5_1x2 xcut143 
transform 1 0 4937 0 1 2431
box 4937 2431 4971 2527
use SUNSAR_cut_M1M4_2x1 xcut144 
transform 1 0 5967 0 1 555
box 5967 555 6059 589
use SUNSAR_cut_M4M5_1x2 xcut145 
transform 1 0 6207 0 1 555
box 6207 555 6241 651
use SUNSAR_cut_M4M5_1x2 xcut146 
transform 1 0 6207 0 1 2431
box 6207 2431 6241 2527
use SUNSAR_cut_M1M3_2x1 xcut147 
transform 1 0 5103 0 1 1259
box 5103 1259 5195 1293
use SUNSAR_cut_M1M3_2x1 xcut148 
transform 1 0 5967 0 1 555
box 5967 555 6059 589
use SUNSAR_cut_M1M4_2x1 xcut149 
transform 1 0 5103 0 1 555
box 5103 555 5195 589
use SUNSAR_cut_M1M4_2x1 xcut150 
transform 1 0 5967 0 1 1259
box 5967 1259 6059 1293
use SUNSAR_cut_M1M3_2x1 xcut151 
transform 1 0 81 0 1 13738
box 81 13738 173 13772
<< labels >>
flabel m3 s 97 9978 131 14354 0 FreeSans 400 0 0 0 D<7>
port 6 nsew signal bidirectional
flabel m3 s 1881 10350 1915 14369 0 FreeSans 400 0 0 0 D<6>
port 7 nsew signal bidirectional
flabel m3 s 2962 10443 2996 14369 0 FreeSans 400 0 0 0 D<5>
port 8 nsew signal bidirectional
flabel m3 s 4401 10536 4435 14369 0 FreeSans 400 0 0 0 D<4>
port 9 nsew signal bidirectional
flabel m3 s 5482 10629 5516 14369 0 FreeSans 400 0 0 0 D<3>
port 10 nsew signal bidirectional
flabel m3 s 6921 10722 6955 14369 0 FreeSans 400 0 0 0 D<2>
port 11 nsew signal bidirectional
flabel m3 s 8002 10815 8036 14369 0 FreeSans 400 0 0 0 D<1>
port 12 nsew signal bidirectional
flabel m1 s 11581 -360 11673 17811 0 FreeSans 400 0 0 0 AVSS
port 19 nsew signal bidirectional
flabel m1 s 11941 -720 12033 18171 0 FreeSans 400 0 0 0 AVDD
port 18 nsew signal bidirectional
flabel m1 s -855 18439 12033 18531 0 FreeSans 400 0 0 0 VREF
port 17 nsew signal bidirectional
flabel m1 s 12105 -826 12139 18531 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 16 nsew signal bidirectional
flabel locali s 9513 16334 9621 16368 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel m3 s 5103 115 5195 149 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel m3 s 5983 115 6075 149 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s 81 15762 189 15796 0 FreeSans 400 0 0 0 CK_SAMPLE
port 15 nsew signal bidirectional
flabel locali s 909 13738 1017 13772 0 FreeSans 400 0 0 0 EN
port 14 nsew signal bidirectional
flabel locali s 5103 1259 5211 1293 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 5103 555 5211 589 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel m3 s 9441 14369 9475 14461 0 FreeSans 400 0 0 0 D<0>
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -961 -932 12139 18531
<< end >>
