magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 68 0 5786 6978
<< m1 >>
rect 914 5282 948 6944
rect 914 5282 948 6944
rect 820 74 854 6944
rect 820 74 854 6944
rect 726 2116 760 6944
rect 726 2116 760 6944
rect 632 3852 666 6944
rect 632 3852 666 6944
rect 538 3546 572 6944
rect 538 3546 572 6944
rect 444 4464 478 6944
rect 444 4464 478 6944
rect 350 2728 384 6944
rect 350 2728 384 6944
rect 256 3034 290 6944
rect 256 3034 290 6944
rect 162 2422 196 6944
rect 162 2422 196 6944
rect 68 3340 102 6944
rect 68 3340 102 6944
rect 1034 1810 1068 1902
rect 1034 1837 1198 1871
rect 1198 0 5748 38
<< m2 >>
rect 948 5309 1034 5347
rect 948 6839 1034 6877
rect 948 5921 1034 5959
rect 948 6533 1034 6571
rect 948 6227 1034 6265
rect 948 5615 1034 5653
rect 854 101 1034 139
rect 854 1631 1034 1669
rect 854 713 1034 751
rect 854 1325 1034 1363
rect 854 1019 1034 1057
rect 854 407 1034 445
rect 760 2143 1034 2181
rect 666 3879 1034 3917
rect 572 3573 1034 3611
rect 572 5103 1034 5141
rect 572 4185 1034 4223
rect 572 4797 1034 4835
rect 478 4491 1034 4529
rect 384 2755 1034 2793
rect 290 3061 1034 3099
rect 196 2449 1034 2487
rect 102 3367 1034 3405
<< locali >>
rect 1034 1810 1068 1902
<< viali >>
rect 1037 1816 1065 1844
rect 1037 1868 1065 1896
<< m3 >>
rect 1198 5208 1236 6978
use SUNSAR_CAP32C_CV XC1 
transform 1 0 1034 0 1 0
box 1034 0 5786 1736
use SUNSAR_CAP32C_CV XC32a<0> 
transform 1 0 1034 0 1 1736
box 1034 1736 5786 3472
use SUNSAR_CAP32C_CV X16ab 
transform 1 0 1034 0 1 3472
box 1034 3472 5786 5208
use SUNSAR_CAP32C_CV XC0 
transform 1 0 1034 0 1 5208
box 1034 5208 5786 6944
use SUNSAR_cut_M1M3_2x1 xcut0 
transform 1 0 1034 0 1 5309
box 1034 5309 1126 5343
use SUNSAR_cut_M2M3_1x2 xcut1 
transform 1 0 914 0 1 5282
box 914 5282 948 5374
use SUNSAR_cut_M1M3_2x1 xcut2 
transform 1 0 1034 0 1 6839
box 1034 6839 1126 6873
use SUNSAR_cut_M2M3_1x2 xcut3 
transform 1 0 914 0 1 6812
box 914 6812 948 6904
use SUNSAR_cut_M1M3_2x1 xcut4 
transform 1 0 1034 0 1 5921
box 1034 5921 1126 5955
use SUNSAR_cut_M2M3_1x2 xcut5 
transform 1 0 914 0 1 5894
box 914 5894 948 5986
use SUNSAR_cut_M1M3_2x1 xcut6 
transform 1 0 1034 0 1 6533
box 1034 6533 1126 6567
use SUNSAR_cut_M2M3_1x2 xcut7 
transform 1 0 914 0 1 6506
box 914 6506 948 6598
use SUNSAR_cut_M1M3_2x1 xcut8 
transform 1 0 1034 0 1 6227
box 1034 6227 1126 6261
use SUNSAR_cut_M2M3_1x2 xcut9 
transform 1 0 914 0 1 6200
box 914 6200 948 6292
use SUNSAR_cut_M1M3_2x1 xcut10 
transform 1 0 1034 0 1 5615
box 1034 5615 1126 5649
use SUNSAR_cut_M2M3_1x2 xcut11 
transform 1 0 914 0 1 5588
box 914 5588 948 5680
use SUNSAR_cut_M1M3_2x1 xcut12 
transform 1 0 1034 0 1 101
box 1034 101 1126 135
use SUNSAR_cut_M2M3_1x2 xcut13 
transform 1 0 820 0 1 74
box 820 74 854 166
use SUNSAR_cut_M1M3_2x1 xcut14 
transform 1 0 1034 0 1 1631
box 1034 1631 1126 1665
use SUNSAR_cut_M2M3_1x2 xcut15 
transform 1 0 820 0 1 1604
box 820 1604 854 1696
use SUNSAR_cut_M1M3_2x1 xcut16 
transform 1 0 1034 0 1 713
box 1034 713 1126 747
use SUNSAR_cut_M2M3_1x2 xcut17 
transform 1 0 820 0 1 686
box 820 686 854 778
use SUNSAR_cut_M1M3_2x1 xcut18 
transform 1 0 1034 0 1 1325
box 1034 1325 1126 1359
use SUNSAR_cut_M2M3_1x2 xcut19 
transform 1 0 820 0 1 1298
box 820 1298 854 1390
use SUNSAR_cut_M1M3_2x1 xcut20 
transform 1 0 1034 0 1 1019
box 1034 1019 1126 1053
use SUNSAR_cut_M2M3_1x2 xcut21 
transform 1 0 820 0 1 992
box 820 992 854 1084
use SUNSAR_cut_M1M3_2x1 xcut22 
transform 1 0 1034 0 1 407
box 1034 407 1126 441
use SUNSAR_cut_M2M3_1x2 xcut23 
transform 1 0 820 0 1 380
box 820 380 854 472
use SUNSAR_cut_M1M3_2x1 xcut24 
transform 1 0 1034 0 1 2143
box 1034 2143 1126 2177
use SUNSAR_cut_M2M3_1x2 xcut25 
transform 1 0 726 0 1 2116
box 726 2116 760 2208
use SUNSAR_cut_M1M3_2x1 xcut26 
transform 1 0 1034 0 1 3879
box 1034 3879 1126 3913
use SUNSAR_cut_M2M3_1x2 xcut27 
transform 1 0 632 0 1 3852
box 632 3852 666 3944
use SUNSAR_cut_M1M3_2x1 xcut28 
transform 1 0 1034 0 1 3573
box 1034 3573 1126 3607
use SUNSAR_cut_M2M3_1x2 xcut29 
transform 1 0 538 0 1 3546
box 538 3546 572 3638
use SUNSAR_cut_M1M3_2x1 xcut30 
transform 1 0 1034 0 1 5103
box 1034 5103 1126 5137
use SUNSAR_cut_M2M3_1x2 xcut31 
transform 1 0 538 0 1 5076
box 538 5076 572 5168
use SUNSAR_cut_M1M3_2x1 xcut32 
transform 1 0 1034 0 1 4185
box 1034 4185 1126 4219
use SUNSAR_cut_M2M3_1x2 xcut33 
transform 1 0 538 0 1 4158
box 538 4158 572 4250
use SUNSAR_cut_M1M3_2x1 xcut34 
transform 1 0 1034 0 1 4797
box 1034 4797 1126 4831
use SUNSAR_cut_M2M3_1x2 xcut35 
transform 1 0 538 0 1 4770
box 538 4770 572 4862
use SUNSAR_cut_M1M3_2x1 xcut36 
transform 1 0 1034 0 1 4491
box 1034 4491 1126 4525
use SUNSAR_cut_M2M3_1x2 xcut37 
transform 1 0 444 0 1 4464
box 444 4464 478 4556
use SUNSAR_cut_M1M3_2x1 xcut38 
transform 1 0 1034 0 1 2755
box 1034 2755 1126 2789
use SUNSAR_cut_M2M3_1x2 xcut39 
transform 1 0 350 0 1 2728
box 350 2728 384 2820
use SUNSAR_cut_M1M3_2x1 xcut40 
transform 1 0 1034 0 1 3061
box 1034 3061 1126 3095
use SUNSAR_cut_M2M3_1x2 xcut41 
transform 1 0 256 0 1 3034
box 256 3034 290 3126
use SUNSAR_cut_M1M3_2x1 xcut42 
transform 1 0 1034 0 1 2449
box 1034 2449 1126 2483
use SUNSAR_cut_M2M3_1x2 xcut43 
transform 1 0 162 0 1 2422
box 162 2422 196 2514
use SUNSAR_cut_M1M3_2x1 xcut44 
transform 1 0 1034 0 1 3367
box 1034 3367 1126 3401
use SUNSAR_cut_M2M3_1x2 xcut45 
transform 1 0 68 0 1 3340
box 68 3340 102 3432
<< labels >>
flabel m1 s 914 5282 948 6944 0 FreeSans 400 0 0 0 CP<9>
port 1 nsew signal bidirectional
flabel m1 s 820 74 854 6944 0 FreeSans 400 0 0 0 CP<8>
port 2 nsew signal bidirectional
flabel m1 s 726 2116 760 6944 0 FreeSans 400 0 0 0 CP<7>
port 3 nsew signal bidirectional
flabel m1 s 632 3852 666 6944 0 FreeSans 400 0 0 0 CP<6>
port 4 nsew signal bidirectional
flabel m1 s 538 3546 572 6944 0 FreeSans 400 0 0 0 CP<5>
port 5 nsew signal bidirectional
flabel m1 s 444 4464 478 6944 0 FreeSans 400 0 0 0 CP<4>
port 6 nsew signal bidirectional
flabel m1 s 350 2728 384 6944 0 FreeSans 400 0 0 0 CP<3>
port 7 nsew signal bidirectional
flabel m1 s 256 3034 290 6944 0 FreeSans 400 0 0 0 CP<2>
port 8 nsew signal bidirectional
flabel m1 s 162 2422 196 6944 0 FreeSans 400 0 0 0 CP<1>
port 9 nsew signal bidirectional
flabel m1 s 68 3340 102 6944 0 FreeSans 400 0 0 0 CP<0>
port 10 nsew signal bidirectional
flabel m1 s 1198 0 5748 38 0 FreeSans 400 0 0 0 AVSS
port 12 nsew signal bidirectional
flabel m3 s 1198 5208 1236 6978 0 FreeSans 400 0 0 0 CTOP
port 11 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 68 0 5786 6978
<< end >>
