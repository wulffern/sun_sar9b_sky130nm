magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 1260 264
<< locali >>
rect 432 203 516 237
rect 516 115 828 149
rect 516 115 550 237
rect 415 115 449 149
rect 162 71 270 105
rect 162 159 270 193
rect 378 203 486 237
rect 1206 66 1314 110
rect -54 66 54 110
<< poly >>
rect 162 79 1098 97
rect 162 167 1098 185
<< m3 >>
rect 774 0 874 264
rect 378 0 478 264
rect 774 0 874 264
rect 378 0 478 264
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 88
box 0 88 630 264
use SUNSAR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNSAR_PCHDL MP1 
transform 1 0 630 0 1 88
box 630 88 1260 264
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 27
box 774 27 874 65
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 203
box 774 203 874 241
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 27
box 378 27 478 65
<< labels >>
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 162 159 270 193 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 378 203 486 237 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 4 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 5 nsew signal bidirectional
flabel m3 s 774 0 874 264 0 FreeSans 400 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel m3 s 378 0 478 264 0 FreeSans 400 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 264
<< end >>
