magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 100 100
<< m1 >>
rect 0 0 92 92
<< v1 >>
rect 6 6 34 34
rect 6 58 34 86
rect 58 6 86 34
rect 58 58 86 86
<< m2 >>
rect 0 0 92 92
<< v2 >>
rect 6 6 34 34
rect 6 58 34 86
rect 58 6 86 34
rect 58 58 86 86
<< m3 >>
rect 0 0 100 100
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 100 100
<< end >>
