magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect -2848 -1848 26216 41790
<< m3 >>
rect 9100 19960 24378 20036
rect 9100 20348 24378 20424
rect 20828 20728 20904 27456
rect 21108 20728 21184 33792
rect 684 20812 760 30968
rect 684 20812 760 30968
rect 4844 21006 4920 30968
rect 5724 21200 5800 30968
rect 1399 21394 1475 30994
rect 4252 21588 4328 30994
rect 4252 21588 4328 30994
rect 6439 21782 6515 30994
rect 6439 21782 6515 30994
rect 9292 21976 9368 30994
rect 9292 21976 9368 30994
rect 11479 22170 11555 30994
rect 11479 22170 11555 30994
rect 14332 22364 14408 30994
rect 14332 22364 14408 30994
rect 16519 22558 16595 30994
rect 16519 22558 16595 30994
rect 1559 22752 1635 32402
rect 4092 22946 4168 32402
rect 6599 23140 6675 32402
rect 1734 23334 1810 33810
rect 3918 23528 3994 33810
rect 6774 23722 6850 33810
rect 8958 23916 9034 33810
rect 11814 24110 11890 33810
rect 13998 24304 14074 33810
rect 16854 24498 16930 33810
rect 1100 25198 1300 40350
rect 4428 25198 4628 40350
rect 6140 25198 6340 40350
rect 9468 25198 9668 40350
rect 11180 25198 11380 40350
rect 14508 25198 14708 40350
rect 16220 25198 16420 40350
rect 19548 25198 19748 40350
rect 21260 25198 21460 40350
rect 9288 -720 9488 5280
rect 13880 -720 14080 5280
rect 1892 25198 2092 41070
rect 3636 25198 3836 41070
rect 6932 25198 7132 41070
rect 8676 25198 8876 41070
rect 11972 25198 12172 41070
rect 13716 25198 13916 41070
rect 17012 25198 17212 41070
rect 18756 25198 18956 41070
rect 22052 25198 22252 41070
rect 8496 -1440 8696 5280
rect 14672 -1440 14872 5280
rect 2468 30008 2668 41790
rect 3060 30008 3260 41790
rect 7508 30008 7708 41790
rect 8100 30008 8300 41790
rect 12548 30008 12748 41790
rect 13140 30008 13340 41790
rect 17588 30008 17788 41790
rect 18180 30008 18380 41790
rect 9934 -1848 10010 3470
rect 13358 -1848 13434 3470
rect 10564 1114 10820 1190
rect 9138 5474 10564 5550
rect 12548 1114 12728 1190
rect 12728 5474 14190 5550
rect 10820 1114 11000 1190
rect 11000 2522 12548 2598
rect 11000 1114 11076 2598
rect 10712 226 10912 302
rect 12456 226 12656 302
rect 19372 30994 19448 31194
<< m2 >>
rect 14152 19454 14228 20036
rect 9100 19454 9176 20424
rect 684 20736 13660 20812
rect 4844 20930 13300 21006
rect 5724 21124 12940 21200
rect 1399 21318 9760 21394
rect 4252 21512 10120 21588
rect 6439 21706 10480 21782
rect 9292 21900 10840 21976
rect 10944 22094 11555 22170
rect 11124 22288 14408 22364
rect 11304 22482 16595 22558
rect 1559 22676 9940 22752
rect 4092 22870 10300 22946
rect 6599 23064 10660 23140
rect 1734 23258 13480 23334
rect 3918 23452 13120 23528
rect 6774 23646 12760 23722
rect 8958 23840 12580 23916
rect 11814 24034 12400 24110
rect 12144 24228 14074 24304
rect 11964 24422 16930 24498
rect 1892 39190 2236 39266
rect 2236 38580 4844 38656
rect 4768 38580 4844 38780
rect 2236 38580 2312 39274
rect 6932 39190 7276 39266
rect 7276 38580 9884 38656
rect 9808 38580 9884 38780
rect 7276 38580 7352 39274
rect 11972 39190 12316 39266
rect 12316 38580 14924 38656
rect 14848 38580 14924 38780
rect 12316 38580 12392 39274
rect 17012 39190 17356 39266
rect 17356 38580 19964 38656
rect 19888 38580 19964 38780
rect 17356 38580 17432 39274
rect 668 35412 20180 35488
rect 592 35412 668 35612
rect 4768 35412 4844 35612
rect 5632 35412 5708 35612
rect 9808 35412 9884 35612
rect 10672 35412 10748 35612
rect 14848 35412 14924 35612
rect 15712 35412 15788 35612
rect 19888 35412 19964 35612
rect 1908 25952 2236 26028
rect 2236 25548 4844 25624
rect 4768 25548 4844 25764
rect 2236 25548 2312 26028
rect 6948 25952 7276 26028
rect 7276 25548 9884 25624
rect 9808 25548 9884 25764
rect 7276 25548 7352 26028
rect 11988 25952 12316 26028
rect 12316 25548 14924 25624
rect 14848 25548 14924 25764
rect 12316 25548 12392 26028
rect 17028 25952 17356 26028
rect 17356 25548 19964 25624
rect 19888 25548 19964 25764
rect 17356 25548 17432 26028
rect 3620 25952 3948 26028
rect 3948 25952 4024 26092
rect 3948 26092 5724 26168
rect 5648 25688 5724 26168
rect 8660 25952 8988 26028
rect 8988 25952 9064 26092
rect 8988 26092 10764 26168
rect 10688 25688 10764 26168
rect 13700 25952 14028 26028
rect 14028 25952 14104 26092
rect 14028 26092 15804 26168
rect 15728 25688 15804 26168
rect 18740 25952 19068 26028
rect 19068 25952 19144 26092
rect 684 27740 20164 27816
rect 608 27448 684 27816
rect 4768 27448 4844 27816
rect 5648 27448 5724 27816
rect 9808 27448 9884 27816
rect 10688 27448 10764 27816
rect 14848 27448 14924 27816
rect 15728 27448 15804 27816
rect 19888 27448 19964 27816
rect 668 28220 20180 28296
rect 592 28220 668 28572
rect 4768 28220 4844 28572
rect 5632 28220 5708 28572
rect 9808 28220 9884 28572
rect 10672 28220 10748 28572
rect 14848 28220 14924 28572
rect 15712 28220 15788 28572
rect 19888 28220 19964 28572
rect 884 29216 2324 29276
rect 2324 29216 3404 29276
rect 2324 29216 7580 29276
rect 2324 29216 8444 29276
rect 2324 29216 12620 29276
rect 2324 29216 13484 29276
rect 2324 29216 17660 29276
rect 2324 29216 18524 29276
rect 20696 30742 21368 30818
rect 20104 27524 20696 27600
rect 20696 27524 20772 30818
rect 20064 27448 20164 27524
rect 20072 28512 20244 28588
rect 20244 31492 22112 31568
rect 20244 28512 20320 31568
rect 22052 31416 22160 31492
rect 22592 38016 22764 38092
rect 20072 36256 22764 36332
rect 22764 36256 22840 38092
rect 18848 39160 20380 39236
rect 20380 38750 20936 38826
rect 20380 38750 20456 39236
rect 22344 38368 22592 38444
rect 19640 37048 22344 37124
rect 22344 37048 22420 38444
rect 10820 2522 10992 2598
rect 10992 1114 12548 1190
rect 10992 1114 11068 2598
rect 668 29216 2540 29276
<< m4 >>
rect 20828 20348 20904 20728
rect 21108 19960 21184 20728
rect 10564 1114 10640 5550
rect 12728 1114 12804 5550
<< m1 >>
rect 13584 19394 13660 20736
rect 13224 19394 13300 20930
rect 12864 19394 12940 21124
rect 9684 19394 9760 21318
rect 10044 19394 10120 21512
rect 10404 19394 10480 21706
rect 10764 19394 10840 21900
rect 10944 19394 11020 22094
rect 11124 19394 11200 22288
rect 11304 19394 11380 22482
rect 9864 19394 9940 22676
rect 10224 19394 10300 22870
rect 10584 19394 10660 23064
rect 13404 19394 13480 23258
rect 13044 19394 13120 23452
rect 12684 19394 12760 23646
rect 12504 19394 12580 23840
rect 12324 19394 12400 24034
rect 12144 19394 12220 24228
rect 11964 19394 12040 24422
rect 9782 -1644 9842 558
rect 13526 -1644 13586 558
rect -2788 38720 668 38780
rect 3620 39160 3956 39220
rect 3956 38600 5708 38660
rect 5648 38600 5708 38780
rect 3956 38600 4016 39228
rect 8660 39160 8996 39220
rect 8996 38600 10748 38660
rect 10688 38600 10748 38780
rect 8996 38600 9056 39228
rect 13700 39160 14036 39220
rect 14036 38600 15788 38660
rect 15728 38600 15788 38780
rect 14036 38600 14096 39228
rect -1924 5474 76 5534
rect -1924 8954 76 9014
rect -1924 12434 76 12494
rect -1924 15914 76 15974
rect 23252 5474 25292 5534
rect 23252 8954 25292 9014
rect 23252 12434 25292 12494
rect 23252 15914 25292 15974
<< locali >>
rect 25092 -720 25292 40350
rect -1924 -720 25292 -520
rect -1924 40150 25292 40350
rect -1924 -720 -1724 40350
rect 25092 -720 25292 40350
rect 25812 -1440 26012 41070
rect -2644 -1440 26012 -1240
rect -2644 40870 26012 41070
rect -2644 -1440 -2444 41070
rect 25812 -1440 26012 41070
rect -2644 41590 26012 41790
rect -2644 41590 26012 41790
rect 26156 -1644 26216 41790
rect -2644 -1644 26216 -1584
rect 26156 -1644 26216 41790
rect -2848 -1848 26216 -1788
rect -2848 -1848 -2788 41790
rect 19532 37048 19748 37108
rect 668 35552 884 35612
rect 2324 29216 2540 29276
rect 10712 2522 10928 2582
rect 10712 1114 10928 1174
use SUNSAR_SARBSSW_CV XB1 
transform -1 0 11684 0 1 0
box 11684 0 24572 5280
use SUNSAR_SARBSSW_CV XB2 
transform 1 0 11684 0 1 0
box 11684 0 24572 5280
use SUNSAR_CDAC7_CV XDAC1 
transform -1 0 11484 0 1 5474
box 11484 5474 22856 19454
use SUNSAR_CDAC7_CV XDAC2 
transform 1 0 11844 0 1 5474
box 11844 5474 23216 19454
use SUNSAR_SARDIGEX4_CV XA0 
transform 1 0 344 0 1 25198
box 344 25198 2864 39630
use SUNSAR_SARDIGEX4_CV XA1 
transform -1 0 5384 0 1 25198
box 5384 25198 7904 39630
use SUNSAR_SARDIGEX4_CV XA2 
transform 1 0 5384 0 1 25198
box 5384 25198 7904 39630
use SUNSAR_SARDIGEX4_CV XA3 
transform -1 0 10424 0 1 25198
box 10424 25198 12944 39630
use SUNSAR_SARDIGEX4_CV XA4 
transform 1 0 10424 0 1 25198
box 10424 25198 12944 39630
use SUNSAR_SARDIGEX4_CV XA5 
transform -1 0 15464 0 1 25198
box 15464 25198 17984 39630
use SUNSAR_SARDIGEX4_CV XA6 
transform 1 0 15464 0 1 25198
box 15464 25198 17984 39630
use SUNSAR_SARDIGEX4_CV XA7 
transform -1 0 20504 0 1 25198
box 20504 25198 23024 39630
use SUNSAR_SARCMPX2_CV XA20 
transform 1 0 20504 0 1 25198
box 20504 25198 23024 39278
use SUNSAR_cut_M3M4_1x2 xcut0 
transform 1 0 14152 0 1 19454
box 14152 19454 14228 19654
use SUNSAR_cut_M3M4_2x1 xcut1 
transform 1 0 14152 0 1 19960
box 14152 19960 14352 20036
use SUNSAR_cut_M3M4_1x2 xcut2 
transform 1 0 9100 0 1 19454
box 9100 19454 9176 19654
use SUNSAR_cut_M3M4_2x1 xcut3 
transform 1 0 9100 0 1 20348
box 9100 20348 9300 20424
use SUNSAR_cut_M2M4_2x1 xcut4 
transform 1 0 20828 0 1 27456
box 20828 27456 21028 27532
use SUNSAR_cut_M4M5_2x1 xcut5 
transform 1 0 20828 0 1 20348
box 20828 20348 21028 20424
use SUNSAR_cut_M4M5_1x2 xcut6 
transform 1 0 20828 0 1 20728
box 20828 20728 20904 20928
use SUNSAR_cut_M3M4_2x1 xcut7 
transform 1 0 20984 0 1 33792
box 20984 33792 21184 33868
use SUNSAR_cut_M2M3_2x1 xcut8 
transform 1 0 20828 0 1 33792
box 20828 33792 21028 33868
use SUNSAR_cut_M4M5_2x1 xcut9 
transform 1 0 21108 0 1 19960
box 21108 19960 21308 20036
use SUNSAR_cut_M4M5_1x2 xcut10 
transform 1 0 21108 0 1 20728
box 21108 20728 21184 20928
use SUNSAR_cut_M3M4_1x2 xcut11 
transform 1 0 684 0 1 20674
box 684 20674 760 20874
use SUNSAR_cut_M2M3_1x2 xcut12 
transform 1 0 13576 0 1 20674
box 13576 20674 13652 20874
use SUNSAR_cut_M3M4_1x2 xcut13 
transform 1 0 4844 0 1 20868
box 4844 20868 4920 21068
use SUNSAR_cut_M2M3_1x2 xcut14 
transform 1 0 13216 0 1 20868
box 13216 20868 13292 21068
use SUNSAR_cut_M3M4_1x2 xcut15 
transform 1 0 5724 0 1 21062
box 5724 21062 5800 21262
use SUNSAR_cut_M2M3_1x2 xcut16 
transform 1 0 12856 0 1 21062
box 12856 21062 12932 21262
use SUNSAR_cut_M3M4_1x2 xcut17 
transform 1 0 1399 0 1 21256
box 1399 21256 1475 21456
use SUNSAR_cut_M2M3_1x2 xcut18 
transform 1 0 9676 0 1 21256
box 9676 21256 9752 21456
use SUNSAR_cut_M3M4_1x2 xcut19 
transform 1 0 4252 0 1 21450
box 4252 21450 4328 21650
use SUNSAR_cut_M2M3_1x2 xcut20 
transform 1 0 10036 0 1 21450
box 10036 21450 10112 21650
use SUNSAR_cut_M3M4_1x2 xcut21 
transform 1 0 6439 0 1 21644
box 6439 21644 6515 21844
use SUNSAR_cut_M2M3_1x2 xcut22 
transform 1 0 10396 0 1 21644
box 10396 21644 10472 21844
use SUNSAR_cut_M3M4_1x2 xcut23 
transform 1 0 9292 0 1 21838
box 9292 21838 9368 22038
use SUNSAR_cut_M2M3_1x2 xcut24 
transform 1 0 10756 0 1 21838
box 10756 21838 10832 22038
use SUNSAR_cut_M3M4_1x2 xcut25 
transform 1 0 11479 0 1 22032
box 11479 22032 11555 22232
use SUNSAR_cut_M2M3_1x2 xcut26 
transform 1 0 10936 0 1 22032
box 10936 22032 11012 22232
use SUNSAR_cut_M3M4_1x2 xcut27 
transform 1 0 14332 0 1 22226
box 14332 22226 14408 22426
use SUNSAR_cut_M2M3_1x2 xcut28 
transform 1 0 11116 0 1 22226
box 11116 22226 11192 22426
use SUNSAR_cut_M3M4_1x2 xcut29 
transform 1 0 16519 0 1 22420
box 16519 22420 16595 22620
use SUNSAR_cut_M2M3_1x2 xcut30 
transform 1 0 11296 0 1 22420
box 11296 22420 11372 22620
use SUNSAR_cut_M3M4_1x2 xcut31 
transform 1 0 1559 0 1 22614
box 1559 22614 1635 22814
use SUNSAR_cut_M2M3_1x2 xcut32 
transform 1 0 9856 0 1 22614
box 9856 22614 9932 22814
use SUNSAR_cut_M3M4_1x2 xcut33 
transform 1 0 4092 0 1 22808
box 4092 22808 4168 23008
use SUNSAR_cut_M2M3_1x2 xcut34 
transform 1 0 10216 0 1 22808
box 10216 22808 10292 23008
use SUNSAR_cut_M3M4_1x2 xcut35 
transform 1 0 6599 0 1 23002
box 6599 23002 6675 23202
use SUNSAR_cut_M2M3_1x2 xcut36 
transform 1 0 10576 0 1 23002
box 10576 23002 10652 23202
use SUNSAR_cut_M3M4_1x2 xcut37 
transform 1 0 1734 0 1 23196
box 1734 23196 1810 23396
use SUNSAR_cut_M2M3_1x2 xcut38 
transform 1 0 13396 0 1 23196
box 13396 23196 13472 23396
use SUNSAR_cut_M3M4_1x2 xcut39 
transform 1 0 3918 0 1 23390
box 3918 23390 3994 23590
use SUNSAR_cut_M2M3_1x2 xcut40 
transform 1 0 13036 0 1 23390
box 13036 23390 13112 23590
use SUNSAR_cut_M3M4_1x2 xcut41 
transform 1 0 6774 0 1 23584
box 6774 23584 6850 23784
use SUNSAR_cut_M2M3_1x2 xcut42 
transform 1 0 12676 0 1 23584
box 12676 23584 12752 23784
use SUNSAR_cut_M3M4_1x2 xcut43 
transform 1 0 8958 0 1 23778
box 8958 23778 9034 23978
use SUNSAR_cut_M2M3_1x2 xcut44 
transform 1 0 12496 0 1 23778
box 12496 23778 12572 23978
use SUNSAR_cut_M3M4_1x2 xcut45 
transform 1 0 11814 0 1 23972
box 11814 23972 11890 24172
use SUNSAR_cut_M2M3_1x2 xcut46 
transform 1 0 12316 0 1 23972
box 12316 23972 12392 24172
use SUNSAR_cut_M3M4_1x2 xcut47 
transform 1 0 13998 0 1 24166
box 13998 24166 14074 24366
use SUNSAR_cut_M2M3_1x2 xcut48 
transform 1 0 12136 0 1 24166
box 12136 24166 12212 24366
use SUNSAR_cut_M3M4_1x2 xcut49 
transform 1 0 16854 0 1 24360
box 16854 24360 16930 24560
use SUNSAR_cut_M2M3_1x2 xcut50 
transform 1 0 11956 0 1 24360
box 11956 24360 12032 24560
use SUNSAR_cut_M1M4_2x2 xcut51 
transform 1 0 1100 0 1 40150
box 1100 40150 1300 40350
use SUNSAR_cut_M1M4_2x2 xcut52 
transform 1 0 4428 0 1 40150
box 4428 40150 4628 40350
use SUNSAR_cut_M1M4_2x2 xcut53 
transform 1 0 6140 0 1 40150
box 6140 40150 6340 40350
use SUNSAR_cut_M1M4_2x2 xcut54 
transform 1 0 9468 0 1 40150
box 9468 40150 9668 40350
use SUNSAR_cut_M1M4_2x2 xcut55 
transform 1 0 11180 0 1 40150
box 11180 40150 11380 40350
use SUNSAR_cut_M1M4_2x2 xcut56 
transform 1 0 14508 0 1 40150
box 14508 40150 14708 40350
use SUNSAR_cut_M1M4_2x2 xcut57 
transform 1 0 16220 0 1 40150
box 16220 40150 16420 40350
use SUNSAR_cut_M1M4_2x2 xcut58 
transform 1 0 19548 0 1 40150
box 19548 40150 19748 40350
use SUNSAR_cut_M1M4_2x2 xcut59 
transform 1 0 21260 0 1 40150
box 21260 40150 21460 40350
use SUNSAR_cut_M1M4_2x2 xcut60 
transform 1 0 9288 0 1 -720
box 9288 -720 9488 -520
use SUNSAR_cut_M1M4_2x2 xcut61 
transform 1 0 13880 0 1 -720
box 13880 -720 14080 -520
use SUNSAR_cut_M1M4_2x2 xcut62 
transform 1 0 1892 0 1 40870
box 1892 40870 2092 41070
use SUNSAR_cut_M1M4_2x2 xcut63 
transform 1 0 3636 0 1 40870
box 3636 40870 3836 41070
use SUNSAR_cut_M1M4_2x2 xcut64 
transform 1 0 6932 0 1 40870
box 6932 40870 7132 41070
use SUNSAR_cut_M1M4_2x2 xcut65 
transform 1 0 8676 0 1 40870
box 8676 40870 8876 41070
use SUNSAR_cut_M1M4_2x2 xcut66 
transform 1 0 11972 0 1 40870
box 11972 40870 12172 41070
use SUNSAR_cut_M1M4_2x2 xcut67 
transform 1 0 13716 0 1 40870
box 13716 40870 13916 41070
use SUNSAR_cut_M1M4_2x2 xcut68 
transform 1 0 17012 0 1 40870
box 17012 40870 17212 41070
use SUNSAR_cut_M1M4_2x2 xcut69 
transform 1 0 18756 0 1 40870
box 18756 40870 18956 41070
use SUNSAR_cut_M1M4_2x2 xcut70 
transform 1 0 22052 0 1 40870
box 22052 40870 22252 41070
use SUNSAR_cut_M1M4_2x2 xcut71 
transform 1 0 8496 0 1 -1440
box 8496 -1440 8696 -1240
use SUNSAR_cut_M1M4_2x2 xcut72 
transform 1 0 14672 0 1 -1440
box 14672 -1440 14872 -1240
use SUNSAR_cut_M1M4_2x2 xcut73 
transform 1 0 2468 0 1 41590
box 2468 41590 2668 41790
use SUNSAR_cut_M1M4_2x2 xcut74 
transform 1 0 3060 0 1 41590
box 3060 41590 3260 41790
use SUNSAR_cut_M1M4_2x2 xcut75 
transform 1 0 7508 0 1 41590
box 7508 41590 7708 41790
use SUNSAR_cut_M1M4_2x2 xcut76 
transform 1 0 8100 0 1 41590
box 8100 41590 8300 41790
use SUNSAR_cut_M1M4_2x2 xcut77 
transform 1 0 12548 0 1 41590
box 12548 41590 12748 41790
use SUNSAR_cut_M1M4_2x2 xcut78 
transform 1 0 13140 0 1 41590
box 13140 41590 13340 41790
use SUNSAR_cut_M1M4_2x2 xcut79 
transform 1 0 17588 0 1 41590
box 17588 41590 17788 41790
use SUNSAR_cut_M1M4_2x2 xcut80 
transform 1 0 18180 0 1 41590
box 18180 41590 18380 41790
use SUNSAR_cut_M1M2_2x1 xcut81 
transform 1 0 9720 0 1 498
box 9720 498 9904 566
use SUNSAR_cut_M1M2_2x1 xcut82 
transform 1 0 9720 0 1 -1644
box 9720 -1644 9904 -1576
use SUNSAR_cut_M1M2_2x1 xcut83 
transform 1 0 13464 0 1 498
box 13464 498 13648 566
use SUNSAR_cut_M1M2_2x1 xcut84 
transform 1 0 13464 0 1 -1644
box 13464 -1644 13648 -1576
use SUNSAR_cut_M1M2_2x1 xcut85 
transform 1 0 668 0 1 38720
box 668 38720 852 38788
use SUNSAR_cut_M1M2_1x2 xcut86 
transform 1 0 -2852 0 1 38658
box -2852 38658 -2784 38842
use SUNSAR_cut_M1M4_2x1 xcut87 
transform 1 0 9872 0 1 -1848
box 9872 -1848 10072 -1772
use SUNSAR_cut_M1M4_2x1 xcut88 
transform 1 0 13296 0 1 -1848
box 13296 -1848 13496 -1772
use SUNSAR_cut_M1M3_2x1 xcut89 
transform 1 0 1892 0 1 39198
box 1892 39198 2092 39274
use SUNSAR_cut_M1M3_2x1 xcut90 
transform 1 0 4844 0 1 38720
box 4844 38720 5044 38796
use SUNSAR_cut_M1M3_2x1 xcut91 
transform 1 0 6932 0 1 39198
box 6932 39198 7132 39274
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 9884 0 1 38720
box 9884 38720 10084 38796
use SUNSAR_cut_M1M3_2x1 xcut93 
transform 1 0 11972 0 1 39198
box 11972 39198 12172 39274
use SUNSAR_cut_M1M3_2x1 xcut94 
transform 1 0 14924 0 1 38720
box 14924 38720 15124 38796
use SUNSAR_cut_M1M3_2x1 xcut95 
transform 1 0 17012 0 1 39198
box 17012 39198 17212 39274
use SUNSAR_cut_M1M3_2x1 xcut96 
transform 1 0 19964 0 1 38720
box 19964 38720 20164 38796
use SUNSAR_cut_M1M3_2x1 xcut97 
transform 1 0 668 0 1 35552
box 668 35552 868 35628
use SUNSAR_cut_M1M3_2x1 xcut98 
transform 1 0 4844 0 1 35552
box 4844 35552 5044 35628
use SUNSAR_cut_M1M3_2x1 xcut99 
transform 1 0 5708 0 1 35552
box 5708 35552 5908 35628
use SUNSAR_cut_M1M3_2x1 xcut100 
transform 1 0 9884 0 1 35552
box 9884 35552 10084 35628
use SUNSAR_cut_M1M3_2x1 xcut101 
transform 1 0 10748 0 1 35552
box 10748 35552 10948 35628
use SUNSAR_cut_M1M3_2x1 xcut102 
transform 1 0 14924 0 1 35552
box 14924 35552 15124 35628
use SUNSAR_cut_M1M3_2x1 xcut103 
transform 1 0 15788 0 1 35552
box 15788 35552 15988 35628
use SUNSAR_cut_M1M3_2x1 xcut104 
transform 1 0 19964 0 1 35552
box 19964 35552 20164 35628
use SUNSAR_cut_M1M2_2x1 xcut105 
transform 1 0 3620 0 1 39160
box 3620 39160 3804 39228
use SUNSAR_cut_M1M2_2x1 xcut106 
transform 1 0 5708 0 1 38720
box 5708 38720 5892 38788
use SUNSAR_cut_M1M2_2x1 xcut107 
transform 1 0 8660 0 1 39160
box 8660 39160 8844 39228
use SUNSAR_cut_M1M2_2x1 xcut108 
transform 1 0 10748 0 1 38720
box 10748 38720 10932 38788
use SUNSAR_cut_M1M2_2x1 xcut109 
transform 1 0 13700 0 1 39160
box 13700 39160 13884 39228
use SUNSAR_cut_M1M2_2x1 xcut110 
transform 1 0 15788 0 1 38720
box 15788 38720 15972 38788
use SUNSAR_cut_M1M3_2x1 xcut111 
transform 1 0 668 0 1 28512
box 668 28512 868 28588
use SUNSAR_cut_M1M3_2x1 xcut112 
transform 1 0 4844 0 1 28512
box 4844 28512 5044 28588
use SUNSAR_cut_M1M3_2x1 xcut113 
transform 1 0 5708 0 1 28512
box 5708 28512 5908 28588
use SUNSAR_cut_M1M3_2x1 xcut114 
transform 1 0 9884 0 1 28512
box 9884 28512 10084 28588
use SUNSAR_cut_M1M3_2x1 xcut115 
transform 1 0 10748 0 1 28512
box 10748 28512 10948 28588
use SUNSAR_cut_M1M3_2x1 xcut116 
transform 1 0 14924 0 1 28512
box 14924 28512 15124 28588
use SUNSAR_cut_M1M3_2x1 xcut117 
transform 1 0 15788 0 1 28512
box 15788 28512 15988 28588
use SUNSAR_cut_M1M3_2x1 xcut118 
transform 1 0 19964 0 1 28512
box 19964 28512 20164 28588
use SUNSAR_cut_M1M3_2x1 xcut119 
transform 1 0 2324 0 1 29216
box 2324 29216 2524 29292
use SUNSAR_cut_M1M3_2x1 xcut120 
transform 1 0 3188 0 1 29216
box 3188 29216 3388 29292
use SUNSAR_cut_M1M3_2x1 xcut121 
transform 1 0 7364 0 1 29216
box 7364 29216 7564 29292
use SUNSAR_cut_M1M3_2x1 xcut122 
transform 1 0 8228 0 1 29216
box 8228 29216 8428 29292
use SUNSAR_cut_M1M3_2x1 xcut123 
transform 1 0 12404 0 1 29216
box 12404 29216 12604 29292
use SUNSAR_cut_M1M3_2x1 xcut124 
transform 1 0 13268 0 1 29216
box 13268 29216 13468 29292
use SUNSAR_cut_M1M3_2x1 xcut125 
transform 1 0 17444 0 1 29216
box 17444 29216 17644 29292
use SUNSAR_cut_M1M3_2x1 xcut126 
transform 1 0 18308 0 1 29216
box 18308 29216 18508 29292
use SUNSAR_cut_M1M3_2x1 xcut127 
transform 1 0 21276 0 1 30750
box 21276 30750 21476 30826
use SUNSAR_cut_M1M3_2x1 xcut128 
transform 1 0 22052 0 1 31416
box 22052 31416 22252 31492
use SUNSAR_cut_M1M3_2x1 xcut129 
transform 1 0 22484 0 1 38016
box 22484 38016 22684 38092
use SUNSAR_cut_M1M3_2x1 xcut130 
transform 1 0 19964 0 1 36256
box 19964 36256 20164 36332
use SUNSAR_cut_M1M3_2x1 xcut131 
transform 1 0 18740 0 1 39160
box 18740 39160 18940 39236
use SUNSAR_cut_M1M3_2x1 xcut132 
transform 1 0 20828 0 1 38758
box 20828 38758 21028 38834
use SUNSAR_cut_M1M3_2x1 xcut133 
transform 1 0 22500 0 1 38368
box 22500 38368 22700 38444
use SUNSAR_cut_M1M3_2x1 xcut134 
transform 1 0 19548 0 1 37048
box 19548 37048 19748 37124
use SUNSAR_cut_M4M5_1x2 xcut135 
transform 1 0 10564 0 1 1114
box 10564 1114 10640 1314
use SUNSAR_cut_M4M5_1x2 xcut136 
transform 1 0 10564 0 1 5350
box 10564 5350 10640 5550
use SUNSAR_cut_M1M4_2x1 xcut137 
transform 1 0 12440 0 1 1114
box 12440 1114 12640 1190
use SUNSAR_cut_M4M5_1x2 xcut138 
transform 1 0 12728 0 1 1114
box 12728 1114 12804 1314
use SUNSAR_cut_M4M5_1x2 xcut139 
transform 1 0 12728 0 1 5350
box 12728 5350 12804 5550
use SUNSAR_cut_M1M3_2x1 xcut140 
transform 1 0 10712 0 1 2522
box 10712 2522 10912 2598
use SUNSAR_cut_M1M3_2x1 xcut141 
transform 1 0 12440 0 1 1114
box 12440 1114 12640 1190
use SUNSAR_cut_M1M4_2x1 xcut142 
transform 1 0 10712 0 1 1114
box 10712 1114 10912 1190
use SUNSAR_cut_M1M4_2x1 xcut143 
transform 1 0 12440 0 1 2522
box 12440 2522 12640 2598
use SUNSAR_cut_M1M3_2x1 xcut144 
transform 1 0 668 0 1 29216
box 668 29216 868 29292
use SUNSAR_cut_M1M2_2x2 xcut145 
transform 1 0 -1924 0 1 5534
box -1924 5534 -1740 5718
use SUNSAR_cut_M1M2_2x2 xcut146 
transform 1 0 -1924 0 1 9014
box -1924 9014 -1740 9198
use SUNSAR_cut_M1M2_2x2 xcut147 
transform 1 0 -1924 0 1 12494
box -1924 12494 -1740 12678
use SUNSAR_cut_M1M2_2x2 xcut148 
transform 1 0 -1924 0 1 15974
box -1924 15974 -1740 16158
use SUNSAR_cut_M1M2_1x2 xcut149 
transform 1 0 25224 0 1 5474
box 25224 5474 25292 5658
use SUNSAR_cut_M1M2_1x2 xcut150 
transform 1 0 25224 0 1 8954
box 25224 8954 25292 9138
use SUNSAR_cut_M1M2_1x2 xcut151 
transform 1 0 25224 0 1 12434
box 25224 12434 25292 12618
use SUNSAR_cut_M1M2_1x2 xcut152 
transform 1 0 25224 0 1 15914
box 25224 15914 25292 16098
<< labels >>
flabel m3 s 684 20812 760 30968 0 FreeSans 400 0 0 0 D<7>
port 6 nsew signal bidirectional
flabel m3 s 4252 21588 4328 30994 0 FreeSans 400 0 0 0 D<6>
port 7 nsew signal bidirectional
flabel m3 s 6439 21782 6515 30994 0 FreeSans 400 0 0 0 D<5>
port 8 nsew signal bidirectional
flabel m3 s 9292 21976 9368 30994 0 FreeSans 400 0 0 0 D<4>
port 9 nsew signal bidirectional
flabel m3 s 11479 22170 11555 30994 0 FreeSans 400 0 0 0 D<3>
port 10 nsew signal bidirectional
flabel m3 s 14332 22364 14408 30994 0 FreeSans 400 0 0 0 D<2>
port 11 nsew signal bidirectional
flabel m3 s 16519 22558 16595 30994 0 FreeSans 400 0 0 0 D<1>
port 12 nsew signal bidirectional
flabel locali s 25092 -720 25292 40350 0 FreeSans 400 0 0 0 AVSS
port 19 nsew signal bidirectional
flabel locali s 25812 -1440 26012 41070 0 FreeSans 400 0 0 0 AVDD
port 18 nsew signal bidirectional
flabel locali s -2644 41590 26012 41790 0 FreeSans 400 0 0 0 VREF
port 17 nsew signal bidirectional
flabel locali s 26156 -1644 26216 41790 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 16 nsew signal bidirectional
flabel locali s 19532 37048 19748 37108 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel m3 s 10712 226 10912 302 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel m3 s 12456 226 12656 302 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s 668 35552 884 35612 0 FreeSans 400 0 0 0 CK_SAMPLE
port 15 nsew signal bidirectional
flabel locali s 2324 29216 2540 29276 0 FreeSans 400 0 0 0 EN
port 14 nsew signal bidirectional
flabel locali s 10712 2522 10928 2582 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 10712 1114 10928 1174 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel m3 s 19372 30994 19448 31194 0 FreeSans 400 0 0 0 D<0>
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -2848 26216 -1848 41790
<< end >>
