magic
tech sky130A
timestamp 1712959200
<< checkpaint >>
rect 0 0 92 34
<< metal1 >>
rect 0 31 92 34
rect 0 3 6 31
rect 34 3 58 31
rect 86 3 92 31
rect 0 0 92 3
<< via1 >>
rect 6 3 34 31
rect 58 3 86 31
<< metal2 >>
rect 0 31 92 34
rect 0 3 6 31
rect 34 3 58 31
rect 86 3 92 31
rect 0 0 92 3
<< properties >>
string FIXED_BBOX 0 0 92 34
<< end >>
