magic
tech sky130B
timestamp 1708692311
<< poly >>
rect 162 167 1098 185
rect 162 79 1098 97
<< locali >>
rect 378 291 828 325
rect 162 247 270 281
rect 990 247 1098 281
rect 378 203 882 237
rect -54 154 54 198
rect 162 159 270 193
rect 415 115 449 149
rect 162 71 270 105
rect 710 61 744 203
rect 1206 154 1314 198
rect 710 27 828 61
<< metal3 >>
rect 378 0 470 352
rect 774 0 866 352
use SUNSAR_NCHDL  MN0
timestamp 1708642800
transform 1 0 0 0 1 88
box -90 -66 630 242
use SUNSAR_NCHDL  MN1
timestamp 1708642800
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNSAR_NCHDL  MN2
timestamp 1708642800
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_PCHDL  MP0
timestamp 1708642800
transform 1 0 630 0 1 88
box 0 -66 720 242
use SUNSAR_PCHDL  MP1
timestamp 1708642800
transform 1 0 630 0 1 176
box 0 -66 720 242
use SUNSAR_PCHDL  MP2
timestamp 1708642800
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1708642800
transform 1 0 774 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1708642800
transform 1 0 774 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut2
timestamp 1708642800
transform 1 0 378 0 1 27
box 0 0 92 34
<< labels >>
flabel locali s 162 159 270 193 0 FreeSans 200 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 990 247 1098 281 0 FreeSans 200 0 0 0 CN
port 3 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 200 0 0 0 C
port 2 nsew signal bidirectional
flabel locali s 162 71 270 105 0 FreeSans 200 0 0 0 RN
port 4 nsew signal bidirectional
flabel locali s 378 291 486 325 0 FreeSans 200 0 0 0 Y
port 5 nsew signal bidirectional
flabel locali s 1206 154 1314 198 0 FreeSans 200 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -54 154 54 198 0 FreeSans 200 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel metal3 s 774 0 866 352 0 FreeSans 200 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel metal3 s 378 0 470 352 0 FreeSans 200 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 352
<< end >>
