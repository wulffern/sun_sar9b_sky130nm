magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect -1077 -932 13175 25991
<< m3 >>
rect 4550 16660 12256 16694
rect 4550 16846 12256 16880
rect 12079 17032 12113 20230
rect 12217 17032 12251 22518
rect -81 17066 -47 21812
rect -81 17066 -47 21812
rect 4519 17159 4553 21812
rect 2439 17252 2473 21812
rect 1999 17345 2033 21812
rect 276 17438 310 21825
rect 4223 17531 4257 21825
rect 4223 17531 4257 21825
rect 5316 17624 5350 21825
rect 5316 17624 5350 21825
rect 6743 17717 6777 21825
rect 6743 17717 6777 21825
rect 7836 17810 7870 21825
rect 7836 17810 7870 21825
rect 9263 17903 9297 21825
rect 9263 17903 9297 21825
rect 2796 17996 2830 21825
rect 2796 17996 2830 21825
rect 1703 18089 1737 21825
rect 1703 18089 1737 21825
rect 2876 18182 2910 22265
rect 4143 18275 4177 22265
rect 1623 18368 1657 22265
rect 356 18461 390 22265
rect 444 18554 478 22705
rect 1536 18647 1570 22705
rect 2964 18740 2998 22705
rect 4056 18833 4090 22705
rect 5484 18926 5518 22705
rect 6576 19019 6610 22705
rect 8004 19112 8038 22705
rect 9096 19205 9130 22705
rect 127 19543 227 25271
rect 1791 19543 1891 25271
rect 2647 19543 2747 25271
rect 4311 19543 4411 25271
rect 5167 19543 5267 25271
rect 6831 19543 6931 25271
rect 7687 19543 7787 25271
rect 9351 19543 9451 25271
rect 10207 19543 10307 25271
rect 11871 19543 11971 25271
rect 4851 -360 4951 2400
rect 7147 -360 7247 2400
rect 523 19543 623 25631
rect 1395 19543 1495 25631
rect 3043 19543 3143 25631
rect 3915 19543 4015 25631
rect 5563 19543 5663 25631
rect 6435 19543 6535 25631
rect 8083 19543 8183 25631
rect 8955 19543 9055 25631
rect 10603 19543 10703 25631
rect 11475 19543 11575 25631
rect 4455 -720 4555 2400
rect 7543 -720 7643 2400
rect 811 21506 911 25991
rect 1107 21506 1207 25991
rect 3331 21506 3431 25991
rect 3627 21506 3727 25991
rect 5851 21506 5951 25991
rect 6147 21506 6247 25991
rect 8371 21506 8471 25991
rect 8667 21506 8767 25991
rect 10891 21506 10991 25991
rect 5176 -932 5210 1471
rect 6888 -932 6922 1471
rect 5397 555 5617 589
rect 4569 2493 5397 2527
rect 6481 555 6667 589
rect 6667 2493 7529 2527
rect 5617 555 5701 589
rect 5701 1259 6481 1293
rect 5701 555 5735 1293
rect 5563 113 5663 151
rect 6435 113 6535 151
rect 10356 21825 10394 21925
<< m2 >>
rect 7510 16415 7544 16698
rect 4550 16415 4584 16884
rect -81 17032 7260 17066
rect 4519 17125 6696 17159
rect 2439 17218 6884 17252
rect 1999 17311 7072 17345
rect 276 17404 4872 17438
rect 4223 17497 5436 17531
rect 5316 17590 5624 17624
rect 5684 17683 6777 17717
rect 5778 17776 7870 17810
rect 5872 17869 9297 17903
rect 2796 17962 5248 17996
rect 1703 18055 5060 18089
rect 2876 18148 5342 18182
rect 4143 18241 5530 18275
rect 1623 18334 5154 18368
rect 356 18427 4966 18461
rect 444 18520 7166 18554
rect 1536 18613 6978 18647
rect 2964 18706 6790 18740
rect 4056 18799 6602 18833
rect 5484 18892 6508 18926
rect 6380 18985 6610 19019
rect 6286 19078 8038 19112
rect 6192 19171 9130 19205
rect 5096 -826 5130 281
rect 6968 -826 7002 281
rect -1043 24454 -89 24488
rect 523 24691 691 24725
rect 691 24390 1999 24424
rect 1965 24390 1999 24488
rect 691 24390 725 24725
rect 3043 24691 3211 24725
rect 3211 24390 4519 24424
rect 4485 24390 4519 24488
rect 3211 24390 3245 24725
rect 5563 24691 5731 24725
rect 5731 24390 7039 24424
rect 7005 24390 7039 24488
rect 5731 24390 5765 24725
rect 8083 24691 8251 24725
rect 8251 24390 9559 24424
rect 9525 24390 9559 24488
rect 8251 24390 8285 24725
rect -89 23158 10099 23192
rect -123 23158 -89 23256
rect 1965 23158 1999 23256
rect 2397 23158 2431 23256
rect 4485 23158 4519 23256
rect 4917 23158 4951 23256
rect 7005 23158 7039 23256
rect 7437 23158 7471 23256
rect 9525 23158 9559 23256
rect 9957 23158 9991 23256
rect 539 19922 691 19956
rect 691 19726 1999 19760
rect 1965 19726 1999 19824
rect 691 19726 725 19956
rect 3059 19922 3211 19956
rect 3211 19726 4519 19760
rect 4485 19726 4519 19824
rect 3211 19726 3245 19956
rect 5579 19922 5731 19956
rect 5731 19726 7039 19760
rect 7005 19726 7039 19824
rect 5731 19726 5765 19956
rect 8099 19922 8251 19956
rect 8251 19726 9559 19760
rect 9525 19726 9559 19824
rect 8251 19726 8285 19956
rect 10619 19922 10771 19956
rect 10771 19922 10805 19956
rect 1387 19922 1539 19956
rect 1539 19922 1573 19986
rect 1539 19986 2447 20020
rect 2413 19790 2447 20020
rect 3907 19922 4059 19956
rect 4059 19922 4093 19986
rect 4059 19986 4967 20020
rect 4933 19790 4967 20020
rect 6427 19922 6579 19956
rect 6579 19922 6613 19986
rect 6579 19986 7487 20020
rect 7453 19790 7487 20020
rect 8947 19922 9099 19956
rect 9099 19922 9133 19986
rect 9099 19986 10007 20020
rect 9973 19790 10007 20020
rect -73 20808 10099 20842
rect -107 20670 -73 20842
rect 1965 20670 1999 20842
rect 2413 20670 2447 20842
rect 4485 20670 4519 20842
rect 4933 20670 4967 20842
rect 7005 20670 7039 20842
rect 7453 20670 7487 20842
rect 9525 20670 9559 20842
rect 9973 20670 10007 20842
rect -89 20884 10099 20918
rect -123 20884 -89 21056
rect 1965 20884 1999 21056
rect 2397 20884 2431 21056
rect 4485 20884 4519 21056
rect 4917 20884 4951 21056
rect 7005 20884 7039 21056
rect 7437 20884 7471 21056
rect 9525 20884 9559 21056
rect 9957 20884 9991 21056
rect 19 21198 739 21232
rect 739 21198 1279 21232
rect 739 21198 3367 21232
rect 739 21198 3799 21232
rect 739 21198 5887 21232
rect 739 21198 6319 21232
rect 739 21198 8407 21232
rect 739 21198 8839 21232
rect 739 21198 10927 21232
rect 11193 21259 11917 21293
rect 10069 20704 11193 20738
rect 11193 20704 11227 21293
rect 10053 20670 10099 20704
rect 11085 21699 11521 21733
rect 10069 21056 11085 21090
rect 11085 21056 11119 21733
rect 10045 21022 10099 21056
rect 11305 23926 11389 23960
rect 10045 23398 11389 23432
rect 11389 23398 11423 23960
rect 11187 24190 11305 24224
rect 10657 24691 11187 24725
rect 11187 24190 11221 24725
rect 5617 1259 5701 1293
rect 5701 555 6481 589
rect 5701 555 5735 1293
rect -89 21198 847 21232
<< m4 >>
rect 12079 16846 12113 17032
rect 12217 16660 12251 17032
rect 5397 555 5431 2527
rect 6667 555 6701 2527
<< m1 >>
rect 7226 16381 7260 17032
rect 6662 16381 6696 17125
rect 6850 16381 6884 17218
rect 7038 16381 7072 17311
rect 4838 16381 4872 17404
rect 5402 16381 5436 17497
rect 5590 16381 5624 17590
rect 5684 16381 5718 17683
rect 5778 16381 5812 17776
rect 5872 16381 5906 17869
rect 5214 16381 5248 17962
rect 5026 16381 5060 18055
rect 5308 16381 5342 18148
rect 5496 16381 5530 18241
rect 5120 16381 5154 18334
rect 4932 16381 4966 18427
rect 7132 16381 7166 18520
rect 6944 16381 6978 18613
rect 6756 16381 6790 18706
rect 6568 16381 6602 18799
rect 6474 16381 6508 18892
rect 6380 16381 6414 18985
rect 6286 16381 6320 19078
rect 6192 16381 6226 19171
rect 12609 -360 12709 25271
rect -611 -360 12709 -260
rect -611 25171 12709 25271
rect -611 -360 -511 25271
rect 12609 -360 12709 25271
rect 12969 -720 13069 25631
rect -971 -720 13069 -620
rect -971 25531 13069 25631
rect -971 -720 -871 25631
rect 12969 -720 13069 25631
rect -971 25891 13069 25991
rect -971 25891 13069 25991
rect 13141 -826 13175 25991
rect -971 -826 13175 -792
rect 13141 -826 13175 25991
rect -1077 -932 13175 -898
rect -1077 -932 -1043 25991
rect 1387 24674 1555 24708
rect 1555 24390 2431 24424
rect 2397 24390 2431 24488
rect 1555 24390 1589 24708
rect 3907 24674 4075 24708
rect 4075 24390 4951 24424
rect 4917 24390 4951 24488
rect 4075 24390 4109 24708
rect 6427 24674 6595 24708
rect 6595 24390 7471 24424
rect 7437 24390 7471 24488
rect 6595 24390 6629 24708
rect 8947 24674 9115 24708
rect 9115 24390 9991 24424
rect 9957 24390 9991 24488
rect 9115 24390 9149 24708
rect 11187 24014 11305 24048
rect 10261 23794 11187 23828
rect 11187 23794 11221 24048
rect -611 2493 38 2527
rect -611 4229 38 4263
rect -611 5965 38 5999
rect -611 7701 38 7735
rect -611 9437 38 9471
rect -611 11173 38 11207
rect -611 12909 38 12943
rect -611 14645 38 14679
rect 12060 2493 12709 2527
rect 12060 4229 12709 4263
rect 12060 5965 12709 5999
rect 12060 7701 12709 7735
rect 12060 9437 12709 9471
rect 12060 11173 12709 11207
rect 12060 12909 12709 12943
rect 12060 14645 12709 14679
<< locali >>
rect 10207 23794 10315 23828
rect -89 23222 19 23256
rect 739 21198 847 21232
rect 5563 1259 5671 1293
rect 5563 555 5671 589
use SUNSAR_SARBSSW_CV XB1 
transform -1 0 6049 0 1 0
box 6049 0 11773 2400
use SUNSAR_SARBSSW_CV XB2 
transform 1 0 6049 0 1 0
box 6049 0 11773 2400
use SUNSAR_CDAC8_CV XDAC1 
transform -1 0 5974 0 1 2493
box 5974 2493 11880 16415
use SUNSAR_CDAC8_CV XDAC2 
transform 1 0 6124 0 1 2493
box 6124 2493 12030 16415
use SUNSAR_SARDIGEX4_CV XA0 
transform 1 0 -251 0 1 19543
box -251 19543 1009 24911
use SUNSAR_SARDIGEX4_CV XA1 
transform -1 0 2269 0 1 19543
box 2269 19543 3529 24911
use SUNSAR_SARDIGEX4_CV XA2 
transform 1 0 2269 0 1 19543
box 2269 19543 3529 24911
use SUNSAR_SARDIGEX4_CV XA3 
transform -1 0 4789 0 1 19543
box 4789 19543 6049 24911
use SUNSAR_SARDIGEX4_CV XA4 
transform 1 0 4789 0 1 19543
box 4789 19543 6049 24911
use SUNSAR_SARDIGEX4_CV XA5 
transform -1 0 7309 0 1 19543
box 7309 19543 8569 24911
use SUNSAR_SARDIGEX4_CV XA6 
transform 1 0 7309 0 1 19543
box 7309 19543 8569 24911
use SUNSAR_SARDIGEX4_CV XA7 
transform -1 0 9829 0 1 19543
box 9829 19543 11089 24911
use SUNSAR_SARDIGEX4_CV XA8 
transform 1 0 9829 0 1 19543
box 9829 19543 11089 24911
use SUNSAR_SARCMPX1_CV XA20 
transform -1 0 12349 0 1 19543
box 12349 19543 13609 24471
use SUNSAR_cut_M3M4_1x2 xcut0 
transform 1 0 7510 0 1 16415
box 7510 16415 7548 16515
use SUNSAR_cut_M3M4_2x1 xcut1 
transform 1 0 7510 0 1 16660
box 7510 16660 7610 16698
use SUNSAR_cut_M3M4_1x2 xcut2 
transform 1 0 4550 0 1 16415
box 4550 16415 4588 16515
use SUNSAR_cut_M3M4_2x1 xcut3 
transform 1 0 4550 0 1 16846
box 4550 16846 4650 16884
use SUNSAR_cut_M2M4_2x1 xcut4 
transform 1 0 12079 0 1 20230
box 12079 20230 12179 20268
use SUNSAR_cut_M4M5_2x1 xcut5 
transform 1 0 12079 0 1 16846
box 12079 16846 12179 16884
use SUNSAR_cut_M4M5_1x2 xcut6 
transform 1 0 12079 0 1 17032
box 12079 17032 12117 17132
use SUNSAR_cut_M3M4_2x1 xcut7 
transform 1 0 12159 0 1 22518
box 12159 22518 12259 22556
use SUNSAR_cut_M2M3_2x1 xcut8 
transform 1 0 12079 0 1 22518
box 12079 22518 12171 22552
use SUNSAR_cut_M4M5_2x1 xcut9 
transform 1 0 12217 0 1 16660
box 12217 16660 12317 16698
use SUNSAR_cut_M4M5_1x2 xcut10 
transform 1 0 12217 0 1 17032
box 12217 17032 12255 17132
use SUNSAR_cut_M3M4_1x2 xcut11 
transform 1 0 -83 0 1 16999
box -83 16999 -45 17099
use SUNSAR_cut_M2M3_1x2 xcut12 
transform 1 0 7226 0 1 17003
box 7226 17003 7260 17095
use SUNSAR_cut_M3M4_1x2 xcut13 
transform 1 0 4517 0 1 17092
box 4517 17092 4555 17192
use SUNSAR_cut_M2M3_1x2 xcut14 
transform 1 0 6662 0 1 17096
box 6662 17096 6696 17188
use SUNSAR_cut_M3M4_1x2 xcut15 
transform 1 0 2437 0 1 17185
box 2437 17185 2475 17285
use SUNSAR_cut_M2M3_1x2 xcut16 
transform 1 0 6850 0 1 17189
box 6850 17189 6884 17281
use SUNSAR_cut_M3M4_1x2 xcut17 
transform 1 0 1997 0 1 17278
box 1997 17278 2035 17378
use SUNSAR_cut_M2M3_1x2 xcut18 
transform 1 0 7038 0 1 17282
box 7038 17282 7072 17374
use SUNSAR_cut_M3M4_1x2 xcut19 
transform 1 0 274 0 1 17371
box 274 17371 312 17471
use SUNSAR_cut_M2M3_1x2 xcut20 
transform 1 0 4838 0 1 17375
box 4838 17375 4872 17467
use SUNSAR_cut_M3M4_1x2 xcut21 
transform 1 0 4221 0 1 17464
box 4221 17464 4259 17564
use SUNSAR_cut_M2M3_1x2 xcut22 
transform 1 0 5402 0 1 17468
box 5402 17468 5436 17560
use SUNSAR_cut_M3M4_1x2 xcut23 
transform 1 0 5314 0 1 17557
box 5314 17557 5352 17657
use SUNSAR_cut_M2M3_1x2 xcut24 
transform 1 0 5590 0 1 17561
box 5590 17561 5624 17653
use SUNSAR_cut_M3M4_1x2 xcut25 
transform 1 0 6741 0 1 17650
box 6741 17650 6779 17750
use SUNSAR_cut_M2M3_1x2 xcut26 
transform 1 0 5684 0 1 17654
box 5684 17654 5718 17746
use SUNSAR_cut_M3M4_1x2 xcut27 
transform 1 0 7834 0 1 17743
box 7834 17743 7872 17843
use SUNSAR_cut_M2M3_1x2 xcut28 
transform 1 0 5778 0 1 17747
box 5778 17747 5812 17839
use SUNSAR_cut_M3M4_1x2 xcut29 
transform 1 0 9261 0 1 17836
box 9261 17836 9299 17936
use SUNSAR_cut_M2M3_1x2 xcut30 
transform 1 0 5872 0 1 17840
box 5872 17840 5906 17932
use SUNSAR_cut_M3M4_1x2 xcut31 
transform 1 0 2794 0 1 17929
box 2794 17929 2832 18029
use SUNSAR_cut_M2M3_1x2 xcut32 
transform 1 0 5214 0 1 17933
box 5214 17933 5248 18025
use SUNSAR_cut_M3M4_1x2 xcut33 
transform 1 0 1701 0 1 18022
box 1701 18022 1739 18122
use SUNSAR_cut_M2M3_1x2 xcut34 
transform 1 0 5026 0 1 18026
box 5026 18026 5060 18118
use SUNSAR_cut_M3M4_1x2 xcut35 
transform 1 0 2874 0 1 18115
box 2874 18115 2912 18215
use SUNSAR_cut_M2M3_1x2 xcut36 
transform 1 0 5308 0 1 18119
box 5308 18119 5342 18211
use SUNSAR_cut_M3M4_1x2 xcut37 
transform 1 0 4141 0 1 18208
box 4141 18208 4179 18308
use SUNSAR_cut_M2M3_1x2 xcut38 
transform 1 0 5496 0 1 18212
box 5496 18212 5530 18304
use SUNSAR_cut_M3M4_1x2 xcut39 
transform 1 0 1621 0 1 18301
box 1621 18301 1659 18401
use SUNSAR_cut_M2M3_1x2 xcut40 
transform 1 0 5120 0 1 18305
box 5120 18305 5154 18397
use SUNSAR_cut_M3M4_1x2 xcut41 
transform 1 0 354 0 1 18394
box 354 18394 392 18494
use SUNSAR_cut_M2M3_1x2 xcut42 
transform 1 0 4932 0 1 18398
box 4932 18398 4966 18490
use SUNSAR_cut_M3M4_1x2 xcut43 
transform 1 0 442 0 1 18487
box 442 18487 480 18587
use SUNSAR_cut_M2M3_1x2 xcut44 
transform 1 0 7132 0 1 18491
box 7132 18491 7166 18583
use SUNSAR_cut_M3M4_1x2 xcut45 
transform 1 0 1534 0 1 18580
box 1534 18580 1572 18680
use SUNSAR_cut_M2M3_1x2 xcut46 
transform 1 0 6944 0 1 18584
box 6944 18584 6978 18676
use SUNSAR_cut_M3M4_1x2 xcut47 
transform 1 0 2962 0 1 18673
box 2962 18673 3000 18773
use SUNSAR_cut_M2M3_1x2 xcut48 
transform 1 0 6756 0 1 18677
box 6756 18677 6790 18769
use SUNSAR_cut_M3M4_1x2 xcut49 
transform 1 0 4054 0 1 18766
box 4054 18766 4092 18866
use SUNSAR_cut_M2M3_1x2 xcut50 
transform 1 0 6568 0 1 18770
box 6568 18770 6602 18862
use SUNSAR_cut_M3M4_1x2 xcut51 
transform 1 0 5482 0 1 18859
box 5482 18859 5520 18959
use SUNSAR_cut_M2M3_1x2 xcut52 
transform 1 0 6474 0 1 18863
box 6474 18863 6508 18955
use SUNSAR_cut_M3M4_1x2 xcut53 
transform 1 0 6574 0 1 18952
box 6574 18952 6612 19052
use SUNSAR_cut_M2M3_1x2 xcut54 
transform 1 0 6380 0 1 18956
box 6380 18956 6414 19048
use SUNSAR_cut_M3M4_1x2 xcut55 
transform 1 0 8002 0 1 19045
box 8002 19045 8040 19145
use SUNSAR_cut_M2M3_1x2 xcut56 
transform 1 0 6286 0 1 19049
box 6286 19049 6320 19141
use SUNSAR_cut_M3M4_1x2 xcut57 
transform 1 0 9094 0 1 19138
box 9094 19138 9132 19238
use SUNSAR_cut_M2M3_1x2 xcut58 
transform 1 0 6192 0 1 19142
box 6192 19142 6226 19234
use SUNSAR_cut_M2M4_2x2 xcut59 
transform 1 0 127 0 1 25171
box 127 25171 227 25271
use SUNSAR_cut_M2M4_2x2 xcut60 
transform 1 0 1791 0 1 25171
box 1791 25171 1891 25271
use SUNSAR_cut_M2M4_2x2 xcut61 
transform 1 0 2647 0 1 25171
box 2647 25171 2747 25271
use SUNSAR_cut_M2M4_2x2 xcut62 
transform 1 0 4311 0 1 25171
box 4311 25171 4411 25271
use SUNSAR_cut_M2M4_2x2 xcut63 
transform 1 0 5167 0 1 25171
box 5167 25171 5267 25271
use SUNSAR_cut_M2M4_2x2 xcut64 
transform 1 0 6831 0 1 25171
box 6831 25171 6931 25271
use SUNSAR_cut_M2M4_2x2 xcut65 
transform 1 0 7687 0 1 25171
box 7687 25171 7787 25271
use SUNSAR_cut_M2M4_2x2 xcut66 
transform 1 0 9351 0 1 25171
box 9351 25171 9451 25271
use SUNSAR_cut_M2M4_2x2 xcut67 
transform 1 0 10207 0 1 25171
box 10207 25171 10307 25271
use SUNSAR_cut_M2M4_2x2 xcut68 
transform 1 0 11871 0 1 25171
box 11871 25171 11971 25271
use SUNSAR_cut_M2M4_2x2 xcut69 
transform 1 0 4851 0 1 -360
box 4851 -360 4951 -260
use SUNSAR_cut_M2M4_2x2 xcut70 
transform 1 0 7147 0 1 -360
box 7147 -360 7247 -260
use SUNSAR_cut_M2M4_2x2 xcut71 
transform 1 0 523 0 1 25531
box 523 25531 623 25631
use SUNSAR_cut_M2M4_2x2 xcut72 
transform 1 0 1395 0 1 25531
box 1395 25531 1495 25631
use SUNSAR_cut_M2M4_2x2 xcut73 
transform 1 0 3043 0 1 25531
box 3043 25531 3143 25631
use SUNSAR_cut_M2M4_2x2 xcut74 
transform 1 0 3915 0 1 25531
box 3915 25531 4015 25631
use SUNSAR_cut_M2M4_2x2 xcut75 
transform 1 0 5563 0 1 25531
box 5563 25531 5663 25631
use SUNSAR_cut_M2M4_2x2 xcut76 
transform 1 0 6435 0 1 25531
box 6435 25531 6535 25631
use SUNSAR_cut_M2M4_2x2 xcut77 
transform 1 0 8083 0 1 25531
box 8083 25531 8183 25631
use SUNSAR_cut_M2M4_2x2 xcut78 
transform 1 0 8955 0 1 25531
box 8955 25531 9055 25631
use SUNSAR_cut_M2M4_2x2 xcut79 
transform 1 0 10603 0 1 25531
box 10603 25531 10703 25631
use SUNSAR_cut_M2M4_2x2 xcut80 
transform 1 0 11475 0 1 25531
box 11475 25531 11575 25631
use SUNSAR_cut_M2M4_2x2 xcut81 
transform 1 0 4455 0 1 -720
box 4455 -720 4555 -620
use SUNSAR_cut_M2M4_2x2 xcut82 
transform 1 0 7543 0 1 -720
box 7543 -720 7643 -620
use SUNSAR_cut_M2M4_2x2 xcut83 
transform 1 0 811 0 1 25891
box 811 25891 911 25991
use SUNSAR_cut_M2M4_2x2 xcut84 
transform 1 0 1107 0 1 25891
box 1107 25891 1207 25991
use SUNSAR_cut_M2M4_2x2 xcut85 
transform 1 0 3331 0 1 25891
box 3331 25891 3431 25991
use SUNSAR_cut_M2M4_2x2 xcut86 
transform 1 0 3627 0 1 25891
box 3627 25891 3727 25991
use SUNSAR_cut_M2M4_2x2 xcut87 
transform 1 0 5851 0 1 25891
box 5851 25891 5951 25991
use SUNSAR_cut_M2M4_2x2 xcut88 
transform 1 0 6147 0 1 25891
box 6147 25891 6247 25991
use SUNSAR_cut_M2M4_2x2 xcut89 
transform 1 0 8371 0 1 25891
box 8371 25891 8471 25991
use SUNSAR_cut_M2M4_2x2 xcut90 
transform 1 0 8667 0 1 25891
box 8667 25891 8767 25991
use SUNSAR_cut_M2M4_2x2 xcut91 
transform 1 0 10891 0 1 25891
box 10891 25891 10991 25991
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 5067 0 1 247
box 5067 247 5159 281
use SUNSAR_cut_M2M3_2x1 xcut93 
transform 1 0 5067 0 1 -826
box 5067 -826 5159 -792
use SUNSAR_cut_M1M3_2x1 xcut94 
transform 1 0 6939 0 1 247
box 6939 247 7031 281
use SUNSAR_cut_M2M3_2x1 xcut95 
transform 1 0 6939 0 1 -826
box 6939 -826 7031 -792
use SUNSAR_cut_M1M3_2x1 xcut96 
transform 1 0 -89 0 1 24454
box -89 24454 3 24488
use SUNSAR_cut_M2M3_1x2 xcut97 
transform 1 0 -1077 0 1 24425
box -1077 24425 -1043 24517
use SUNSAR_cut_M2M4_2x1 xcut98 
transform 1 0 5143 0 1 -932
box 5143 -932 5243 -894
use SUNSAR_cut_M2M4_2x1 xcut99 
transform 1 0 6855 0 1 -932
box 6855 -932 6955 -894
use SUNSAR_cut_M1M3_2x1 xcut100 
transform 1 0 523 0 1 24691
box 523 24691 615 24725
use SUNSAR_cut_M1M3_2x1 xcut101 
transform 1 0 1999 0 1 24454
box 1999 24454 2091 24488
use SUNSAR_cut_M1M3_2x1 xcut102 
transform 1 0 3043 0 1 24691
box 3043 24691 3135 24725
use SUNSAR_cut_M1M3_2x1 xcut103 
transform 1 0 4519 0 1 24454
box 4519 24454 4611 24488
use SUNSAR_cut_M1M3_2x1 xcut104 
transform 1 0 5563 0 1 24691
box 5563 24691 5655 24725
use SUNSAR_cut_M1M3_2x1 xcut105 
transform 1 0 7039 0 1 24454
box 7039 24454 7131 24488
use SUNSAR_cut_M1M3_2x1 xcut106 
transform 1 0 8083 0 1 24691
box 8083 24691 8175 24725
use SUNSAR_cut_M1M3_2x1 xcut107 
transform 1 0 9559 0 1 24454
box 9559 24454 9651 24488
use SUNSAR_cut_M1M3_2x1 xcut108 
transform 1 0 -89 0 1 23222
box -89 23222 3 23256
use SUNSAR_cut_M1M3_2x1 xcut109 
transform 1 0 1999 0 1 23222
box 1999 23222 2091 23256
use SUNSAR_cut_M1M3_2x1 xcut110 
transform 1 0 2431 0 1 23222
box 2431 23222 2523 23256
use SUNSAR_cut_M1M3_2x1 xcut111 
transform 1 0 4519 0 1 23222
box 4519 23222 4611 23256
use SUNSAR_cut_M1M3_2x1 xcut112 
transform 1 0 4951 0 1 23222
box 4951 23222 5043 23256
use SUNSAR_cut_M1M3_2x1 xcut113 
transform 1 0 7039 0 1 23222
box 7039 23222 7131 23256
use SUNSAR_cut_M1M3_2x1 xcut114 
transform 1 0 7471 0 1 23222
box 7471 23222 7563 23256
use SUNSAR_cut_M1M3_2x1 xcut115 
transform 1 0 9559 0 1 23222
box 9559 23222 9651 23256
use SUNSAR_cut_M1M3_2x1 xcut116 
transform 1 0 9991 0 1 23222
box 9991 23222 10083 23256
use SUNSAR_cut_M1M2_2x1 xcut117 
transform 1 0 1387 0 1 24674
box 1387 24674 1479 24708
use SUNSAR_cut_M1M2_2x1 xcut118 
transform 1 0 2431 0 1 24454
box 2431 24454 2523 24488
use SUNSAR_cut_M1M2_2x1 xcut119 
transform 1 0 3907 0 1 24674
box 3907 24674 3999 24708
use SUNSAR_cut_M1M2_2x1 xcut120 
transform 1 0 4951 0 1 24454
box 4951 24454 5043 24488
use SUNSAR_cut_M1M2_2x1 xcut121 
transform 1 0 6427 0 1 24674
box 6427 24674 6519 24708
use SUNSAR_cut_M1M2_2x1 xcut122 
transform 1 0 7471 0 1 24454
box 7471 24454 7563 24488
use SUNSAR_cut_M1M2_2x1 xcut123 
transform 1 0 8947 0 1 24674
box 8947 24674 9039 24708
use SUNSAR_cut_M1M2_2x1 xcut124 
transform 1 0 9991 0 1 24454
box 9991 24454 10083 24488
use SUNSAR_cut_M1M3_2x1 xcut125 
transform 1 0 -89 0 1 21022
box -89 21022 3 21056
use SUNSAR_cut_M1M3_2x1 xcut126 
transform 1 0 1999 0 1 21022
box 1999 21022 2091 21056
use SUNSAR_cut_M1M3_2x1 xcut127 
transform 1 0 2431 0 1 21022
box 2431 21022 2523 21056
use SUNSAR_cut_M1M3_2x1 xcut128 
transform 1 0 4519 0 1 21022
box 4519 21022 4611 21056
use SUNSAR_cut_M1M3_2x1 xcut129 
transform 1 0 4951 0 1 21022
box 4951 21022 5043 21056
use SUNSAR_cut_M1M3_2x1 xcut130 
transform 1 0 7039 0 1 21022
box 7039 21022 7131 21056
use SUNSAR_cut_M1M3_2x1 xcut131 
transform 1 0 7471 0 1 21022
box 7471 21022 7563 21056
use SUNSAR_cut_M1M3_2x1 xcut132 
transform 1 0 9559 0 1 21022
box 9559 21022 9651 21056
use SUNSAR_cut_M1M3_2x1 xcut133 
transform 1 0 9991 0 1 21022
box 9991 21022 10083 21056
use SUNSAR_cut_M1M3_2x1 xcut134 
transform 1 0 739 0 1 21198
box 739 21198 831 21232
use SUNSAR_cut_M1M3_2x1 xcut135 
transform 1 0 1171 0 1 21198
box 1171 21198 1263 21232
use SUNSAR_cut_M1M3_2x1 xcut136 
transform 1 0 3259 0 1 21198
box 3259 21198 3351 21232
use SUNSAR_cut_M1M3_2x1 xcut137 
transform 1 0 3691 0 1 21198
box 3691 21198 3783 21232
use SUNSAR_cut_M1M3_2x1 xcut138 
transform 1 0 5779 0 1 21198
box 5779 21198 5871 21232
use SUNSAR_cut_M1M3_2x1 xcut139 
transform 1 0 6211 0 1 21198
box 6211 21198 6303 21232
use SUNSAR_cut_M1M3_2x1 xcut140 
transform 1 0 8299 0 1 21198
box 8299 21198 8391 21232
use SUNSAR_cut_M1M3_2x1 xcut141 
transform 1 0 8731 0 1 21198
box 8731 21198 8823 21232
use SUNSAR_cut_M1M3_2x1 xcut142 
transform 1 0 10819 0 1 21198
box 10819 21198 10911 21232
use SUNSAR_cut_M1M3_2x1 xcut143 
transform 1 0 11879 0 1 21259
box 11879 21259 11971 21293
use SUNSAR_cut_M1M3_2x1 xcut144 
transform 1 0 11483 0 1 21699
box 11483 21699 11575 21733
use SUNSAR_cut_M1M3_2x1 xcut145 
transform 1 0 11251 0 1 23926
box 11251 23926 11343 23960
use SUNSAR_cut_M1M3_2x1 xcut146 
transform 1 0 9991 0 1 23398
box 9991 23398 10083 23432
use SUNSAR_cut_M1M3_2x1 xcut147 
transform 1 0 11267 0 1 24190
box 11267 24190 11359 24224
use SUNSAR_cut_M1M3_2x1 xcut148 
transform 1 0 10619 0 1 24691
box 10619 24691 10711 24725
use SUNSAR_cut_M1M2_2x1 xcut149 
transform 1 0 11267 0 1 24014
box 11267 24014 11359 24048
use SUNSAR_cut_M1M2_2x1 xcut150 
transform 1 0 10223 0 1 23794
box 10223 23794 10315 23828
use SUNSAR_cut_M4M5_1x2 xcut151 
transform 1 0 5397 0 1 555
box 5397 555 5435 655
use SUNSAR_cut_M4M5_1x2 xcut152 
transform 1 0 5397 0 1 2427
box 5397 2427 5435 2527
use SUNSAR_cut_M1M4_2x1 xcut153 
transform 1 0 6427 0 1 555
box 6427 555 6527 593
use SUNSAR_cut_M4M5_1x2 xcut154 
transform 1 0 6667 0 1 555
box 6667 555 6705 655
use SUNSAR_cut_M4M5_1x2 xcut155 
transform 1 0 6667 0 1 2427
box 6667 2427 6705 2527
use SUNSAR_cut_M1M3_2x1 xcut156 
transform 1 0 5563 0 1 1259
box 5563 1259 5655 1293
use SUNSAR_cut_M1M3_2x1 xcut157 
transform 1 0 6427 0 1 555
box 6427 555 6519 589
use SUNSAR_cut_M1M4_2x1 xcut158 
transform 1 0 5563 0 1 555
box 5563 555 5663 593
use SUNSAR_cut_M1M4_2x1 xcut159 
transform 1 0 6427 0 1 1259
box 6427 1259 6527 1297
use SUNSAR_cut_M1M3_2x1 xcut160 
transform 1 0 -89 0 1 21198
box -89 21198 3 21232
<< labels >>
flabel m3 s -81 17066 -47 21812 0 FreeSans 400 0 0 0 D<8>
port 6 nsew signal bidirectional
flabel m3 s 4223 17531 4257 21825 0 FreeSans 400 0 0 0 D<5>
port 9 nsew signal bidirectional
flabel m3 s 5316 17624 5350 21825 0 FreeSans 400 0 0 0 D<4>
port 10 nsew signal bidirectional
flabel m3 s 6743 17717 6777 21825 0 FreeSans 400 0 0 0 D<3>
port 11 nsew signal bidirectional
flabel m3 s 7836 17810 7870 21825 0 FreeSans 400 0 0 0 D<2>
port 12 nsew signal bidirectional
flabel m3 s 9263 17903 9297 21825 0 FreeSans 400 0 0 0 D<1>
port 13 nsew signal bidirectional
flabel m3 s 2796 17996 2830 21825 0 FreeSans 400 0 0 0 D<6>
port 8 nsew signal bidirectional
flabel m3 s 1703 18089 1737 21825 0 FreeSans 400 0 0 0 D<7>
port 7 nsew signal bidirectional
flabel m1 s 12609 -360 12709 25271 0 FreeSans 400 0 0 0 AVSS
port 20 nsew signal bidirectional
flabel m1 s 12969 -720 13069 25631 0 FreeSans 400 0 0 0 AVDD
port 19 nsew signal bidirectional
flabel m1 s -971 25891 13069 25991 0 FreeSans 400 0 0 0 VREF
port 18 nsew signal bidirectional
flabel m1 s 13141 -826 13175 25991 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew signal bidirectional
flabel locali s 10207 23794 10315 23828 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel m3 s 5563 113 5663 151 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel m3 s 6435 113 6535 151 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s -89 23222 19 23256 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew signal bidirectional
flabel locali s 739 21198 847 21232 0 FreeSans 400 0 0 0 EN
port 15 nsew signal bidirectional
flabel locali s 5563 1259 5671 1293 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 5563 555 5671 589 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel m3 s 10356 21825 10394 21925 0 FreeSans 400 0 0 0 D<0>
port 14 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -1077 -932 13175 25991
<< end >>
