magic
tech sky130B
magscale 1 2
timestamp 1708642800
<< checkpaint >>
rect 0 0 7272 960
<< m1 >>
rect 108 -40 7236 40
rect 7164 40 7236 120
rect 108 120 7092 200
rect 7164 120 7236 200
rect 108 200 180 280
rect 7164 200 7236 280
rect 108 280 180 360
rect 252 280 7236 360
rect 108 360 180 440
rect 7164 360 7236 440
rect 108 440 7092 520
rect 7164 440 7236 520
rect 108 520 180 600
rect 7164 520 7236 600
rect 108 600 180 680
rect 252 600 7236 680
rect 108 680 180 760
rect 108 760 7236 840
<< m2 >>
rect 108 -40 7236 40
rect 7164 40 7236 120
rect 108 120 7092 200
rect 7164 120 7236 200
rect 108 200 180 280
rect 7164 200 7236 280
rect 108 280 180 360
rect 252 280 7236 360
rect 108 360 180 440
rect 7164 360 7236 440
rect 108 440 7092 520
rect 7164 440 7236 520
rect 108 520 180 600
rect 7164 520 7236 600
rect 108 600 180 680
rect 252 600 7236 680
rect 108 680 180 760
rect 108 760 7236 840
<< locali >>
rect 108 -40 7236 40
rect 7164 40 7236 120
rect 108 120 7092 200
rect 7164 120 7236 200
rect 108 200 180 280
rect 7164 200 7236 280
rect 108 280 180 360
rect 252 280 7236 360
rect 108 360 180 440
rect 7164 360 7236 440
rect 108 440 7092 520
rect 7164 440 7236 520
rect 108 520 180 600
rect 7164 520 7236 600
rect 108 600 180 680
rect 252 600 7236 680
rect 108 680 180 760
rect 108 760 7236 840
<< v1 >>
rect 6876 -32 6948 -24
rect 6876 -24 6948 -16
rect 6876 -16 6948 -8
rect 6876 -8 6948 0
rect 6876 0 6948 8
rect 6876 8 6948 16
rect 6876 16 6948 24
rect 6876 24 6948 32
rect 6948 -32 7020 -24
rect 6948 -24 7020 -16
rect 6948 -16 7020 -8
rect 6948 -8 7020 0
rect 6948 0 7020 8
rect 6948 8 7020 16
rect 6948 16 7020 24
rect 6948 24 7020 32
rect 7020 -32 7092 -24
rect 7020 -24 7092 -16
rect 7020 -16 7092 -8
rect 7020 -8 7092 0
rect 7020 0 7092 8
rect 7020 8 7092 16
rect 7020 16 7092 24
rect 7020 24 7092 32
rect 324 128 396 136
rect 324 136 396 144
rect 324 144 396 152
rect 324 152 396 160
rect 324 160 396 168
rect 324 168 396 176
rect 324 176 396 184
rect 324 184 396 192
rect 396 128 468 136
rect 396 136 468 144
rect 396 144 468 152
rect 396 152 468 160
rect 396 160 468 168
rect 396 168 468 176
rect 396 176 468 184
rect 396 184 468 192
rect 468 128 540 136
rect 468 136 540 144
rect 468 144 540 152
rect 468 152 540 160
rect 468 160 540 168
rect 468 168 540 176
rect 468 176 540 184
rect 468 184 540 192
rect 6876 288 6948 296
rect 6876 296 6948 304
rect 6876 304 6948 312
rect 6876 312 6948 320
rect 6876 320 6948 328
rect 6876 328 6948 336
rect 6876 336 6948 344
rect 6876 344 6948 352
rect 6948 288 7020 296
rect 6948 296 7020 304
rect 6948 304 7020 312
rect 6948 312 7020 320
rect 6948 320 7020 328
rect 6948 328 7020 336
rect 6948 336 7020 344
rect 6948 344 7020 352
rect 7020 288 7092 296
rect 7020 296 7092 304
rect 7020 304 7092 312
rect 7020 312 7092 320
rect 7020 320 7092 328
rect 7020 328 7092 336
rect 7020 336 7092 344
rect 7020 344 7092 352
rect 324 448 396 456
rect 324 456 396 464
rect 324 464 396 472
rect 324 472 396 480
rect 324 480 396 488
rect 324 488 396 496
rect 324 496 396 504
rect 324 504 396 512
rect 396 448 468 456
rect 396 456 468 464
rect 396 464 468 472
rect 396 472 468 480
rect 396 480 468 488
rect 396 488 468 496
rect 396 496 468 504
rect 396 504 468 512
rect 468 448 540 456
rect 468 456 540 464
rect 468 464 540 472
rect 468 472 540 480
rect 468 480 540 488
rect 468 488 540 496
rect 468 496 540 504
rect 468 504 540 512
rect 6876 608 6948 616
rect 6876 616 6948 624
rect 6876 624 6948 632
rect 6876 632 6948 640
rect 6876 640 6948 648
rect 6876 648 6948 656
rect 6876 656 6948 664
rect 6876 664 6948 672
rect 6948 608 7020 616
rect 6948 616 7020 624
rect 6948 624 7020 632
rect 6948 632 7020 640
rect 6948 640 7020 648
rect 6948 648 7020 656
rect 6948 656 7020 664
rect 6948 664 7020 672
rect 7020 608 7092 616
rect 7020 616 7092 624
rect 7020 624 7092 632
rect 7020 632 7092 640
rect 7020 640 7092 648
rect 7020 648 7092 656
rect 7020 656 7092 664
rect 7020 664 7092 672
rect 324 768 396 776
rect 324 776 396 784
rect 324 784 396 792
rect 324 792 396 800
rect 324 800 396 808
rect 324 808 396 816
rect 324 816 396 824
rect 324 824 396 832
rect 396 768 468 776
rect 396 776 468 784
rect 396 784 468 792
rect 396 792 468 800
rect 396 800 468 808
rect 396 808 468 816
rect 396 816 468 824
rect 396 824 468 832
rect 468 768 540 776
rect 468 776 540 784
rect 468 784 540 792
rect 468 792 540 800
rect 468 800 540 808
rect 468 808 540 816
rect 468 816 540 824
rect 468 824 540 832
<< v2 >>
rect 6876 -32 6948 -24
rect 6876 -24 6948 -16
rect 6876 -16 6948 -8
rect 6876 -8 6948 0
rect 6876 0 6948 8
rect 6876 8 6948 16
rect 6876 16 6948 24
rect 6876 24 6948 32
rect 6948 -32 7020 -24
rect 6948 -24 7020 -16
rect 6948 -16 7020 -8
rect 6948 -8 7020 0
rect 6948 0 7020 8
rect 6948 8 7020 16
rect 6948 16 7020 24
rect 6948 24 7020 32
rect 7020 -32 7092 -24
rect 7020 -24 7092 -16
rect 7020 -16 7092 -8
rect 7020 -8 7092 0
rect 7020 0 7092 8
rect 7020 8 7092 16
rect 7020 16 7092 24
rect 7020 24 7092 32
rect 324 128 396 136
rect 324 136 396 144
rect 324 144 396 152
rect 324 152 396 160
rect 324 160 396 168
rect 324 168 396 176
rect 324 176 396 184
rect 324 184 396 192
rect 396 128 468 136
rect 396 136 468 144
rect 396 144 468 152
rect 396 152 468 160
rect 396 160 468 168
rect 396 168 468 176
rect 396 176 468 184
rect 396 184 468 192
rect 468 128 540 136
rect 468 136 540 144
rect 468 144 540 152
rect 468 152 540 160
rect 468 160 540 168
rect 468 168 540 176
rect 468 176 540 184
rect 468 184 540 192
rect 6876 288 6948 296
rect 6876 296 6948 304
rect 6876 304 6948 312
rect 6876 312 6948 320
rect 6876 320 6948 328
rect 6876 328 6948 336
rect 6876 336 6948 344
rect 6876 344 6948 352
rect 6948 288 7020 296
rect 6948 296 7020 304
rect 6948 304 7020 312
rect 6948 312 7020 320
rect 6948 320 7020 328
rect 6948 328 7020 336
rect 6948 336 7020 344
rect 6948 344 7020 352
rect 7020 288 7092 296
rect 7020 296 7092 304
rect 7020 304 7092 312
rect 7020 312 7092 320
rect 7020 320 7092 328
rect 7020 328 7092 336
rect 7020 336 7092 344
rect 7020 344 7092 352
rect 324 448 396 456
rect 324 456 396 464
rect 324 464 396 472
rect 324 472 396 480
rect 324 480 396 488
rect 324 488 396 496
rect 324 496 396 504
rect 324 504 396 512
rect 396 448 468 456
rect 396 456 468 464
rect 396 464 468 472
rect 396 472 468 480
rect 396 480 468 488
rect 396 488 468 496
rect 396 496 468 504
rect 396 504 468 512
rect 468 448 540 456
rect 468 456 540 464
rect 468 464 540 472
rect 468 472 540 480
rect 468 480 540 488
rect 468 488 540 496
rect 468 496 540 504
rect 468 504 540 512
rect 6876 608 6948 616
rect 6876 616 6948 624
rect 6876 624 6948 632
rect 6876 632 6948 640
rect 6876 640 6948 648
rect 6876 648 6948 656
rect 6876 656 6948 664
rect 6876 664 6948 672
rect 6948 608 7020 616
rect 6948 616 7020 624
rect 6948 624 7020 632
rect 6948 632 7020 640
rect 6948 640 7020 648
rect 6948 648 7020 656
rect 6948 656 7020 664
rect 6948 664 7020 672
rect 7020 608 7092 616
rect 7020 616 7092 624
rect 7020 624 7092 632
rect 7020 632 7092 640
rect 7020 640 7092 648
rect 7020 648 7092 656
rect 7020 656 7092 664
rect 7020 664 7092 672
rect 324 768 396 776
rect 324 776 396 784
rect 324 784 396 792
rect 324 792 396 800
rect 324 800 396 808
rect 324 808 396 816
rect 324 816 396 824
rect 324 824 396 832
rect 396 768 468 776
rect 396 776 468 784
rect 396 784 468 792
rect 396 792 468 800
rect 396 800 468 808
rect 396 808 468 816
rect 396 816 468 824
rect 396 824 468 832
rect 468 768 540 776
rect 468 776 540 784
rect 468 784 540 792
rect 468 792 540 800
rect 468 800 540 808
rect 468 808 540 816
rect 468 816 540 824
rect 468 824 540 832
<< viali >>
rect 6876 -32 6948 -24
rect 6876 -24 6948 -16
rect 6876 -16 6948 -8
rect 6876 -8 6948 0
rect 6876 0 6948 8
rect 6876 8 6948 16
rect 6876 16 6948 24
rect 6876 24 6948 32
rect 6948 -32 7020 -24
rect 6948 -24 7020 -16
rect 6948 -16 7020 -8
rect 6948 -8 7020 0
rect 6948 0 7020 8
rect 6948 8 7020 16
rect 6948 16 7020 24
rect 6948 24 7020 32
rect 7020 -32 7092 -24
rect 7020 -24 7092 -16
rect 7020 -16 7092 -8
rect 7020 -8 7092 0
rect 7020 0 7092 8
rect 7020 8 7092 16
rect 7020 16 7092 24
rect 7020 24 7092 32
rect 324 128 396 136
rect 324 136 396 144
rect 324 144 396 152
rect 324 152 396 160
rect 324 160 396 168
rect 324 168 396 176
rect 324 176 396 184
rect 324 184 396 192
rect 396 128 468 136
rect 396 136 468 144
rect 396 144 468 152
rect 396 152 468 160
rect 396 160 468 168
rect 396 168 468 176
rect 396 176 468 184
rect 396 184 468 192
rect 468 128 540 136
rect 468 136 540 144
rect 468 144 540 152
rect 468 152 540 160
rect 468 160 540 168
rect 468 168 540 176
rect 468 176 540 184
rect 468 184 540 192
rect 6876 288 6948 296
rect 6876 296 6948 304
rect 6876 304 6948 312
rect 6876 312 6948 320
rect 6876 320 6948 328
rect 6876 328 6948 336
rect 6876 336 6948 344
rect 6876 344 6948 352
rect 6948 288 7020 296
rect 6948 296 7020 304
rect 6948 304 7020 312
rect 6948 312 7020 320
rect 6948 320 7020 328
rect 6948 328 7020 336
rect 6948 336 7020 344
rect 6948 344 7020 352
rect 7020 288 7092 296
rect 7020 296 7092 304
rect 7020 304 7092 312
rect 7020 312 7092 320
rect 7020 320 7092 328
rect 7020 328 7092 336
rect 7020 336 7092 344
rect 7020 344 7092 352
rect 324 448 396 456
rect 324 456 396 464
rect 324 464 396 472
rect 324 472 396 480
rect 324 480 396 488
rect 324 488 396 496
rect 324 496 396 504
rect 324 504 396 512
rect 396 448 468 456
rect 396 456 468 464
rect 396 464 468 472
rect 396 472 468 480
rect 396 480 468 488
rect 396 488 468 496
rect 396 496 468 504
rect 396 504 468 512
rect 468 448 540 456
rect 468 456 540 464
rect 468 464 540 472
rect 468 472 540 480
rect 468 480 540 488
rect 468 488 540 496
rect 468 496 540 504
rect 468 504 540 512
rect 6876 608 6948 616
rect 6876 616 6948 624
rect 6876 624 6948 632
rect 6876 632 6948 640
rect 6876 640 6948 648
rect 6876 648 6948 656
rect 6876 656 6948 664
rect 6876 664 6948 672
rect 6948 608 7020 616
rect 6948 616 7020 624
rect 6948 624 7020 632
rect 6948 632 7020 640
rect 6948 640 7020 648
rect 6948 648 7020 656
rect 6948 656 7020 664
rect 6948 664 7020 672
rect 7020 608 7092 616
rect 7020 616 7092 624
rect 7020 624 7092 632
rect 7020 632 7092 640
rect 7020 640 7092 648
rect 7020 648 7092 656
rect 7020 656 7092 664
rect 7020 664 7092 672
rect 324 768 396 776
rect 324 776 396 784
rect 324 784 396 792
rect 324 792 396 800
rect 324 800 396 808
rect 324 808 396 816
rect 324 816 396 824
rect 324 824 396 832
rect 396 768 468 776
rect 396 776 468 784
rect 396 784 468 792
rect 396 792 468 800
rect 396 800 468 808
rect 396 808 468 816
rect 396 816 468 824
rect 396 824 468 832
rect 468 768 540 776
rect 468 776 540 784
rect 468 784 540 792
rect 468 792 540 800
rect 468 800 540 808
rect 468 808 540 816
rect 468 816 540 824
rect 468 824 540 832
<< m3 >>
rect 108 -40 7236 40
rect 108 -40 7236 40
rect 7164 40 7236 120
rect 108 120 6876 200
rect 6948 120 7092 200
rect 7164 120 7236 200
rect 108 200 180 280
rect 7164 200 7236 280
rect 108 280 180 360
rect 252 280 324 360
rect 396 280 7236 360
rect 108 360 180 440
rect 7164 360 7236 440
rect 108 440 7092 520
rect 7164 440 7236 520
rect 108 520 180 600
rect 7164 520 7236 600
rect 108 600 180 680
rect 252 600 7236 680
rect 108 680 180 760
rect 108 760 7236 840
rect 108 760 7236 840
<< rm3 >>
rect 6876 120 6948 200
rect 324 280 396 360
<< v3 >>
rect 6876 -32 6948 -24
rect 6876 -24 6948 -16
rect 6876 -16 6948 -8
rect 6876 -8 6948 0
rect 6876 0 6948 8
rect 6876 8 6948 16
rect 6876 16 6948 24
rect 6876 24 6948 32
rect 6948 -32 7020 -24
rect 6948 -24 7020 -16
rect 6948 -16 7020 -8
rect 6948 -8 7020 0
rect 6948 0 7020 8
rect 6948 8 7020 16
rect 6948 16 7020 24
rect 6948 24 7020 32
rect 7020 -32 7092 -24
rect 7020 -24 7092 -16
rect 7020 -16 7092 -8
rect 7020 -8 7092 0
rect 7020 0 7092 8
rect 7020 8 7092 16
rect 7020 16 7092 24
rect 7020 24 7092 32
rect 324 128 396 136
rect 324 136 396 144
rect 324 144 396 152
rect 324 152 396 160
rect 324 160 396 168
rect 324 168 396 176
rect 324 176 396 184
rect 324 184 396 192
rect 396 128 468 136
rect 396 136 468 144
rect 396 144 468 152
rect 396 152 468 160
rect 396 160 468 168
rect 396 168 468 176
rect 396 176 468 184
rect 396 184 468 192
rect 468 128 540 136
rect 468 136 540 144
rect 468 144 540 152
rect 468 152 540 160
rect 468 160 540 168
rect 468 168 540 176
rect 468 176 540 184
rect 468 184 540 192
rect 6876 288 6948 296
rect 6876 296 6948 304
rect 6876 304 6948 312
rect 6876 312 6948 320
rect 6876 320 6948 328
rect 6876 328 6948 336
rect 6876 336 6948 344
rect 6876 344 6948 352
rect 6948 288 7020 296
rect 6948 296 7020 304
rect 6948 304 7020 312
rect 6948 312 7020 320
rect 6948 320 7020 328
rect 6948 328 7020 336
rect 6948 336 7020 344
rect 6948 344 7020 352
rect 7020 288 7092 296
rect 7020 296 7092 304
rect 7020 304 7092 312
rect 7020 312 7092 320
rect 7020 320 7092 328
rect 7020 328 7092 336
rect 7020 336 7092 344
rect 7020 344 7092 352
rect 324 448 396 456
rect 324 456 396 464
rect 324 464 396 472
rect 324 472 396 480
rect 324 480 396 488
rect 324 488 396 496
rect 324 496 396 504
rect 324 504 396 512
rect 396 448 468 456
rect 396 456 468 464
rect 396 464 468 472
rect 396 472 468 480
rect 396 480 468 488
rect 396 488 468 496
rect 396 496 468 504
rect 396 504 468 512
rect 468 448 540 456
rect 468 456 540 464
rect 468 464 540 472
rect 468 472 540 480
rect 468 480 540 488
rect 468 488 540 496
rect 468 496 540 504
rect 468 504 540 512
rect 6876 608 6948 616
rect 6876 616 6948 624
rect 6876 624 6948 632
rect 6876 632 6948 640
rect 6876 640 6948 648
rect 6876 648 6948 656
rect 6876 656 6948 664
rect 6876 664 6948 672
rect 6948 608 7020 616
rect 6948 616 7020 624
rect 6948 624 7020 632
rect 6948 632 7020 640
rect 6948 640 7020 648
rect 6948 648 7020 656
rect 6948 656 7020 664
rect 6948 664 7020 672
rect 7020 608 7092 616
rect 7020 616 7092 624
rect 7020 624 7092 632
rect 7020 632 7092 640
rect 7020 640 7092 648
rect 7020 648 7092 656
rect 7020 656 7092 664
rect 7020 664 7092 672
rect 324 768 396 776
rect 324 776 396 784
rect 324 784 396 792
rect 324 792 396 800
rect 324 800 396 808
rect 324 808 396 816
rect 324 816 396 824
rect 324 824 396 832
rect 396 768 468 776
rect 396 776 468 784
rect 396 784 468 792
rect 396 792 468 800
rect 396 800 468 808
rect 396 808 468 816
rect 396 816 468 824
rect 396 824 468 832
rect 468 768 540 776
rect 468 776 540 784
rect 468 784 540 792
rect 468 792 540 800
rect 468 800 540 808
rect 468 808 540 816
rect 468 816 540 824
rect 468 824 540 832
<< m4 >>
rect 108 -40 7236 40
rect 7164 40 7236 120
rect 108 120 7092 200
rect 7164 120 7236 200
rect 108 200 180 280
rect 7164 200 7236 280
rect 108 280 180 360
rect 252 280 7236 360
rect 108 360 180 440
rect 7164 360 7236 440
rect 108 440 7092 520
rect 7164 440 7236 520
rect 108 520 180 600
rect 7164 520 7236 600
rect 108 600 180 680
rect 252 600 7236 680
rect 108 680 180 760
rect 108 760 7236 840
<< labels >>
flabel m3 s 108 -40 7236 40 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 108 760 7236 840 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 7272 960
<< end >>
