magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 17 4752 1753
<< m3 >>
rect 164 0 202 1770
rect 164 0 202 1770
rect 234 70 272 1700
rect 304 0 342 1770
rect 374 70 412 1700
rect 444 0 482 1770
rect 514 70 552 1700
rect 584 0 622 1770
rect 654 70 692 1700
rect 724 0 762 1770
rect 794 70 832 1700
rect 864 0 902 1770
rect 934 70 972 1700
rect 1004 0 1042 1770
rect 1074 70 1112 1700
rect 1144 0 1182 1770
rect 1214 70 1252 1700
rect 1284 0 1322 1770
rect 1354 70 1392 1700
rect 1424 0 1462 1770
rect 1494 70 1532 1700
rect 1564 0 1602 1770
rect 1634 70 1672 1700
rect 1704 0 1742 1770
rect 1774 70 1812 1700
rect 1844 0 1882 1770
rect 1914 70 1952 1700
rect 1984 0 2022 1770
rect 2054 70 2092 1700
rect 2124 0 2162 1770
rect 2194 70 2232 1700
rect 2264 0 2302 1770
rect 2334 70 2372 1700
rect 2404 0 2442 1770
rect 2474 70 2512 1700
rect 2544 0 2582 1770
rect 2614 70 2652 1700
rect 2684 0 2722 1770
rect 2754 70 2792 1700
rect 2824 0 2862 1770
rect 2894 70 2932 1700
rect 2964 0 3002 1770
rect 3034 70 3072 1700
rect 3104 0 3142 1770
rect 3174 70 3212 1700
rect 3244 0 3282 1770
rect 3314 70 3352 1700
rect 3384 0 3422 1770
rect 3454 70 3492 1700
rect 3524 0 3562 1770
rect 3594 70 3632 1700
rect 3664 0 3702 1770
rect 3734 70 3772 1700
rect 3804 0 3842 1770
rect 3874 70 3912 1700
rect 3944 0 3982 1770
rect 4014 70 4052 1700
rect 4084 0 4122 1770
rect 4154 70 4192 1700
rect 4224 0 4262 1770
rect 4294 70 4332 1700
rect 4364 0 4402 1770
rect 4434 70 4472 1700
rect 4504 0 4542 1770
rect 4574 70 4612 1700
rect 4714 0 4752 1770
rect 4644 0 4682 1770
rect 164 0 4644 38
rect 164 1732 4644 1770
<< m1 >>
rect 164 0 4714 38
rect 1214 200 1252 1770
rect 3594 0 3632 1570
rect 1354 0 1392 652
rect 1354 812 1392 1770
rect 3454 0 3492 652
rect 3454 812 3492 1770
rect 1074 0 1112 1264
rect 1074 1424 1112 1770
rect 1494 0 1532 1264
rect 1494 1424 1532 1770
rect 3314 0 3352 1264
rect 3314 1424 3352 1770
rect 3734 0 3772 1264
rect 3734 1424 3772 1770
rect 794 0 832 958
rect 794 1118 832 1770
rect 934 0 972 958
rect 934 1118 972 1770
rect 1634 0 1672 958
rect 1634 1118 1672 1770
rect 1774 0 1812 958
rect 1774 1118 1812 1770
rect 3034 0 3072 958
rect 3034 1118 3072 1770
rect 3174 0 3212 958
rect 3174 1118 3212 1770
rect 3874 0 3912 958
rect 3874 1118 3912 1770
rect 4014 0 4052 958
rect 4014 1118 4052 1770
rect 234 0 272 346
rect 234 506 272 1770
rect 374 0 412 346
rect 374 506 412 1770
rect 514 0 552 346
rect 514 506 552 1770
rect 654 0 692 346
rect 654 506 692 1770
rect 1914 0 1952 346
rect 1914 506 1952 1770
rect 2054 0 2092 346
rect 2054 506 2092 1770
rect 2194 0 2232 346
rect 2194 506 2232 1770
rect 2334 0 2372 346
rect 2334 506 2372 1770
rect 2474 0 2512 346
rect 2474 506 2512 1770
rect 2614 0 2652 346
rect 2614 506 2652 1770
rect 2754 0 2792 346
rect 2754 506 2792 1770
rect 2894 0 2932 346
rect 2894 506 2932 1770
rect 4154 0 4192 346
rect 4154 506 4192 1770
rect 4294 0 4332 346
rect 4294 506 4332 1770
rect 4434 0 4472 346
rect 4434 506 4472 1770
rect 4574 0 4612 346
rect 4574 506 4612 1770
rect 164 0 202 1732
rect 304 0 342 1732
rect 444 0 482 1732
rect 584 0 622 1732
rect 724 0 762 1732
rect 864 0 902 1732
rect 1004 0 1042 1732
rect 1144 0 1182 1732
rect 1284 0 1322 1732
rect 1424 0 1462 1732
rect 1564 0 1602 1732
rect 1704 0 1742 1732
rect 1844 0 1882 1732
rect 1984 0 2022 1732
rect 2124 0 2162 1732
rect 2264 0 2302 1732
rect 2404 0 2442 1732
rect 2544 0 2582 1732
rect 2684 0 2722 1732
rect 2824 0 2862 1732
rect 2964 0 3002 1732
rect 3104 0 3142 1732
rect 3244 0 3282 1732
rect 3384 0 3422 1732
rect 3524 0 3562 1732
rect 3664 0 3702 1732
rect 3804 0 3842 1732
rect 3944 0 3982 1732
rect 4084 0 4122 1732
rect 4224 0 4262 1732
rect 4364 0 4402 1732
rect 4504 0 4542 1732
rect 4714 0 4752 1770
rect 4644 0 4682 1770
rect 164 0 4714 38
rect 164 1732 4714 1770
<< locali >>
rect 0 101 100 139
rect 0 1631 100 1669
rect 0 713 100 751
rect 0 1325 100 1363
rect 0 1019 100 1057
rect 0 407 100 445
rect 168 407 4644 445
rect 168 101 4644 139
rect 168 1631 4644 1669
rect 168 713 4644 751
rect 168 1325 4644 1363
rect 168 1019 4644 1057
<< m2 >>
rect 4714 0 4752 1770
use SUNSAR_RM1 XRES1A 
transform 1 0 100 0 1 101
box 100 101 168 135
use SUNSAR_RM1 XRES1B 
transform 1 0 100 0 1 1631
box 100 1631 168 1665
use SUNSAR_RM1 XRES2 
transform 1 0 100 0 1 713
box 100 713 168 747
use SUNSAR_RM1 XRES4 
transform 1 0 100 0 1 1325
box 100 1325 168 1359
use SUNSAR_RM1 XRES8 
transform 1 0 100 0 1 1019
box 100 1019 168 1053
use SUNSAR_RM1 XRES16 
transform 1 0 100 0 1 407
box 100 407 168 441
use SUNSAR_cut_M2M4_1x2 xcut0 
transform 1 0 4714 0 1 785
box 4714 785 4752 885
use SUNSAR_cut_M1M4_1x2 xcut1 
transform 1 0 1214 0 1 70
box 1214 70 1252 170
use SUNSAR_cut_M1M4_1x2 xcut2 
transform 1 0 3594 0 1 1600
box 3594 1600 3632 1700
use SUNSAR_cut_M1M4_1x2 xcut3 
transform 1 0 1354 0 1 682
box 1354 682 1392 782
use SUNSAR_cut_M1M4_1x2 xcut4 
transform 1 0 3454 0 1 682
box 3454 682 3492 782
use SUNSAR_cut_M1M4_1x2 xcut5 
transform 1 0 1074 0 1 1294
box 1074 1294 1112 1394
use SUNSAR_cut_M1M4_1x2 xcut6 
transform 1 0 1494 0 1 1294
box 1494 1294 1532 1394
use SUNSAR_cut_M1M4_1x2 xcut7 
transform 1 0 3314 0 1 1294
box 3314 1294 3352 1394
use SUNSAR_cut_M1M4_1x2 xcut8 
transform 1 0 3734 0 1 1294
box 3734 1294 3772 1394
use SUNSAR_cut_M1M4_1x2 xcut9 
transform 1 0 794 0 1 988
box 794 988 832 1088
use SUNSAR_cut_M1M4_1x2 xcut10 
transform 1 0 934 0 1 988
box 934 988 972 1088
use SUNSAR_cut_M1M4_1x2 xcut11 
transform 1 0 1634 0 1 988
box 1634 988 1672 1088
use SUNSAR_cut_M1M4_1x2 xcut12 
transform 1 0 1774 0 1 988
box 1774 988 1812 1088
use SUNSAR_cut_M1M4_1x2 xcut13 
transform 1 0 3034 0 1 988
box 3034 988 3072 1088
use SUNSAR_cut_M1M4_1x2 xcut14 
transform 1 0 3174 0 1 988
box 3174 988 3212 1088
use SUNSAR_cut_M1M4_1x2 xcut15 
transform 1 0 3874 0 1 988
box 3874 988 3912 1088
use SUNSAR_cut_M1M4_1x2 xcut16 
transform 1 0 4014 0 1 988
box 4014 988 4052 1088
use SUNSAR_cut_M1M4_1x2 xcut17 
transform 1 0 234 0 1 376
box 234 376 272 476
use SUNSAR_cut_M1M4_1x2 xcut18 
transform 1 0 374 0 1 376
box 374 376 412 476
use SUNSAR_cut_M1M4_1x2 xcut19 
transform 1 0 514 0 1 376
box 514 376 552 476
use SUNSAR_cut_M1M4_1x2 xcut20 
transform 1 0 654 0 1 376
box 654 376 692 476
use SUNSAR_cut_M1M4_1x2 xcut21 
transform 1 0 1914 0 1 376
box 1914 376 1952 476
use SUNSAR_cut_M1M4_1x2 xcut22 
transform 1 0 2054 0 1 376
box 2054 376 2092 476
use SUNSAR_cut_M1M4_1x2 xcut23 
transform 1 0 2194 0 1 376
box 2194 376 2232 476
use SUNSAR_cut_M1M4_1x2 xcut24 
transform 1 0 2334 0 1 376
box 2334 376 2372 476
use SUNSAR_cut_M1M4_1x2 xcut25 
transform 1 0 2474 0 1 376
box 2474 376 2512 476
use SUNSAR_cut_M1M4_1x2 xcut26 
transform 1 0 2614 0 1 376
box 2614 376 2652 476
use SUNSAR_cut_M1M4_1x2 xcut27 
transform 1 0 2754 0 1 376
box 2754 376 2792 476
use SUNSAR_cut_M1M4_1x2 xcut28 
transform 1 0 2894 0 1 376
box 2894 376 2932 476
use SUNSAR_cut_M1M4_1x2 xcut29 
transform 1 0 4154 0 1 376
box 4154 376 4192 476
use SUNSAR_cut_M1M4_1x2 xcut30 
transform 1 0 4294 0 1 376
box 4294 376 4332 476
use SUNSAR_cut_M1M4_1x2 xcut31 
transform 1 0 4434 0 1 376
box 4434 376 4472 476
use SUNSAR_cut_M1M4_1x2 xcut32 
transform 1 0 4574 0 1 376
box 4574 376 4612 476
<< labels >>
flabel m3 s 164 0 202 1770 0 FreeSans 400 0 0 0 CTOP
port 7 nsew signal bidirectional
flabel m1 s 164 0 4714 38 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
flabel locali s 0 101 100 139 0 FreeSans 400 0 0 0 C1A
port 1 nsew signal bidirectional
flabel locali s 0 1631 100 1669 0 FreeSans 400 0 0 0 C1B
port 2 nsew signal bidirectional
flabel locali s 0 713 100 751 0 FreeSans 400 0 0 0 C2
port 3 nsew signal bidirectional
flabel locali s 0 1325 100 1363 0 FreeSans 400 0 0 0 C4
port 4 nsew signal bidirectional
flabel locali s 0 1019 100 1057 0 FreeSans 400 0 0 0 C8
port 5 nsew signal bidirectional
flabel locali s 0 407 100 445 0 FreeSans 400 0 0 0 C16
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 17 4752 1753
<< end >>
