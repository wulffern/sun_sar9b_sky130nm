* NGSPICE file created from SUNSAR_SAR9B_CV.ext - technology: sky130B

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0>
+ EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
*.subckt SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4>
*+ D<3> D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
R0 XDAC1.XC128a<1>.XRES16.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X0 XB1.XA4.MN0.G CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X1 AVDD XA4.XA1.XA1.MN0.S XA4.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X2 AVSS XA8.XA3.MN0.G D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X3 XA5.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA6.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X4 XA1.XA10.MN0.G XA1.XA9.MN1.G XA1.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X5 XA0.XA12.MN0.D XA0.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X6 AVDD XA1.XA9.MN1.G XA1.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X7 VREF XA6.XA4.MN0.D XA6.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X8 VREF XA4.XA4.MN0.G XA4.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X9 XA2.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R1 XDAC1.XC64b<1>.XRES1B.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X10 XA5.XA10.MN0.D XA5.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X11 AVSS CK_SAMPLE XA1.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X12 VREF XA6.XA4.MN0.G XA6.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X13 AVDD XA1.XA6.MP0.G XA1.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X14 VREF XA4.XA3.MN0.G D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X15 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X16 XA8.XA9.MN1.G CK_SAMPLE XA8.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X17 XA5.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R2 XA0.XA6.MP0.G XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X18 VREF XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X19 XA20.XA2.MN1.D SARP XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X20 XA20.XA3a.MN0.G XA20.XA3.MN6.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X21 XA6.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X22 XA4.XA9.MN1.G D<4> XA4.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X23 AVSS XA2.XA4.MN0.D XA2.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R3 XDAC1.XC128b<2>.XRES1B.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X24 XA8.XA11.MN1.G XA7.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X25 XA5.XA10.MN0.G XA5.XA9.MN1.G XA5.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X26 XA5.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA5.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X27 XA8.XA11.MN1.G XA7.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X28 XA6.XA4.MN0.D XA6.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X29 AVDD XA20.XA9.MN0.D XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X30 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=227 pd=1.22k as=0.616 ps=3.3 w=1.08 l=0.18
X31 AVSS XA2.XA4.MN0.G XA2.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R4 XDAC1.XC32a<0>.XRES16.B D<6> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X32 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=150 pd=802 as=0.616 ps=3.3 w=1.08 l=0.18
X33 AVSS XA8.XA11.MN1.G XA8.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X34 AVSS CK_SAMPLE XA5.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X35 AVSS XA20.XA3.MN6.D XA20.XA2a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X36 AVDD XA20.XA3.MN6.D XA20.XA2a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X37 VREF XA0.XA1.XA5.MN2.D D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X38 XA20.XA1.MN0.D XA20.XA10.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X39 XA0.XA9.MN0.D XA0.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X40 AVSS XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R5 XDAC1.X16ab.XRES1B.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X41 AVDD XA20.XA10.MN1.D XA20.XA1.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R6 D<8> XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X42 XA8.XA4.MN0.G EN XA8.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X43 XA8.XA7.MN0.D XA8.XA7.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X44 XA20.XA3.MN0.D SARP XA20.XA2.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X45 AVDD XA20.XA3.MN6.D XA20.XA3a.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X46 XA0.XA1.XA4.MP1.D EN XA0.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X47 XA4.XA12.MN0.G XA4.XA11.MN1.G XA4.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X48 VREF XA5.XA4.MN0.D XA5.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X49 XA2.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X50 XA8.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA8.XA7.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X51 XA0.XA6.MP2.G D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X52 SARN XB2.XA4.MN1.D SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X53 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=7.39 ps=39.6 w=1.08 l=0.18
X54 XA6.XA10.MN0.D XA6.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X55 XA2.XA4.MN0.D XA2.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X56 AVDD XB1.XA4.MN0.G XB1.XA3.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X57 AVDD EN XA0.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X58 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X59 XA4.XA7.MN0.D XA5.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X60 VREF XA5.XA3.MN0.G D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X61 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X62 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X63 XA8.XA12.MN0.G XA8.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R7 XDAC1.XC1.XRES1B.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X64 D<8> XA0.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X65 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X66 XA6.XA6.MP2.D D<2> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X67 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X68 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X69 XA7.XA9.MN0.D XA7.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X70 XA7.XA10.MN0.G XA7.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X71 XA3.XA1.XA5.MN2.D XA3.XA1.XA5.MN2.G XA3.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X72 XA3.XA1.XA5.MN2.D EN XA3.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X73 XA0.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X74 XA4.XA11.MP0.D XA4.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X75 XA3.XA4.MN0.D XA3.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R8 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X76 XA3.XA1.XA2.MN0.D XA4.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X77 XA3.XA4.MN0.D XA3.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X78 XA3.XA1.XA2.MN0.D XA4.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X79 AVDD XA6.XA9.MN1.G XA6.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X80 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X81 XA2.XA10.MN0.D XA2.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X82 XA5.XA6.MP0.G XA5.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X83 XA8.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA8.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X84 D<5> XA3.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X85 D<5> XA3.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X86 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=7.39 ps=39.6 w=1.08 l=0.18
X87 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X88 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X89 AVDD XA6.XA6.MP0.G XA6.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X90 XA2.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X91 XA3.XA1.XA5.MN1.D XA3.XA1.XA2.MN0.D XA3.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X92 XA20.XA3.MN1.D SARN XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X93 XA3.XA1.XA5.MP1.D EN XA3.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X94 XA20.XA3.MN1.D XA20.XA9.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X95 XA6.XA4.MN0.G XA6.XA1.XA5.MN2.G XA6.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X96 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X97 XA6.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X98 AVDD XA3.XA1.XA1.MN0.S XA3.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X99 XA0.XA8.MN0.D XA0.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X100 VREF XA8.XA4.MN0.D XA8.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X101 XA2.XA10.MN0.G XA2.XA9.MN1.G XA2.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X102 VREF XA3.XA4.MN0.G XA3.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X103 AVSS XA3.XA4.MN0.G XA3.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X104 XA0.XA6.MP0.G XA0.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X105 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X106 VREF XA8.XA3.MN0.G D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X107 VREF XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X108 AVSS CK_SAMPLE XA2.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X109 AVSS XA3.XA3.MN0.G D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R9 XA0.XA6.MP0.G XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X110 VREF XA3.XA3.MN0.G D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X111 XB2.XA4.MN0.G CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X112 XA2.XA1.XA4.MP1.D EN XA2.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X113 XA6.XA11.MN1.G XA5.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X114 XA4.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X115 D<6> XA2.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X116 AVDD EN XA2.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X117 XA3.XA9.MN1.G CK_SAMPLE XA3.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X118 XA3.XA9.MN1.G D<5> XA3.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X119 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X120 AVSS XA20.XA2a.MN0.D XA6.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X121 XA8.XA6.MP0.G XA8.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X122 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R10 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R11 XDAC1.XC0.XRES2.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R12 D<8> XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X123 XA2.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X124 AVSS XA4.XA4.MN0.D XA4.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R13 XA2.XA6.MP0.G XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X125 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X126 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X127 AVSS XA3.XA11.MN1.G XA3.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X128 AVSS XA6.XA4.MN0.D XA6.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X129 XA3.XA12.MN0.G XA3.XA11.MN1.G XA3.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X130 AVSS XA4.XA4.MN0.G XA4.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X131 XA5.XA10.MN0.G XA5.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X132 XA1.XA1.XA5.MN2.D XA0.XA7.MN0.G XA1.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X133 XA3.XA7.MN0.D XA4.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X134 AVSS XA6.XA3.MN0.G D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X135 AVSS XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X136 XA1.XA1.XA5.MN2.D EN XA1.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X137 XA3.XA7.MN0.D XA4.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R14 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R15 XDAC1.XC64b<1>.XRES8.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X138 XA1.XA4.MN0.D XA1.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X139 XA1.XA4.MN0.D XA1.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R16 XB1.XCAPB1.XCAPB4.B m3_7544_1364# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X140 XA1.XA1.XA2.MN0.D XA2.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X141 XA1.XA1.XA2.MN0.D XA2.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X142 XA4.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R17 XB1.XCAPB1.XCAPB4.B m3_7544_4532# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R18 XB2.XCAPB1.XCAPB4.A m3_26048_3300# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X143 XA20.XA12.MN0.G XA8.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X144 XA2.XA8.MN0.D XA2.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X145 D<7> XA1.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X146 XA3.XA12.MN0.G XA3.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X147 XA0.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X148 XA4.XA4.MN0.D XA4.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X149 D<7> XA1.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X150 XA3.XA11.MP0.D XA3.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X151 XA2.XA6.MP0.G XA2.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X152 XA1.XA1.XA5.MN1.D XA1.XA1.XA2.MN0.D XA1.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X153 D<8> XA0.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X154 XA1.XA1.XA5.MP1.D EN XA1.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X155 XA6.XA6.MP0.G XA6.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X156 XA5.XA1.XA5.MN2.D XA5.XA1.XA5.MN2.G XA5.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X157 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X158 AVDD XA1.XA1.XA1.MN0.S XA1.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X159 XA5.XA4.MN0.D XA5.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X160 AVSS XA1.XA4.MN0.G XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R19 D<8> XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X161 XA5.XA1.XA2.MN0.D XA6.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X162 AVSS XA0.XA4.MN0.D XA0.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X163 VREF XA1.XA4.MN0.G XA1.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X164 XA4.XA10.MN0.D XA4.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X165 XA7.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X166 AVSS XA1.XA3.MN0.G D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X167 D<3> XA5.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R20 m3_16472_1364# XB2.XCAPB1.XCAPB4.B sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X168 XB1.XA4.MN0.D XB1.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X169 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X170 XA7.XA6.MP0.D XA7.XA6.MP0.G XA7.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X171 AVSS XA0.XA4.MN0.G XA0.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X172 VREF XA1.XA3.MN0.G D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R21 XDAC1.XC64b<1>.XRES1A.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R22 m3_16472_4532# XB2.XCAPB1.XCAPB4.B sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X173 XA4.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X174 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X175 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X176 XA5.XA1.XA5.MN1.D XA5.XA1.XA2.MN0.D XA5.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X177 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X178 XA8.XA10.MN0.G XA8.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X179 AVSS XA0.XA1.XA5.MN2.D D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X180 AVSS XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X181 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X182 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X183 XA1.XA9.MN1.G CK_SAMPLE XA1.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X184 XA1.XA9.MN1.G D<7> XA1.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X185 XA0.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X186 XA7.XA11.MN1.G XA6.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X187 XA4.XA10.MN0.G XA4.XA9.MN1.G XA4.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X188 AVSS XA7.XA4.MN0.D XA7.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X189 VREF XA7.XA4.MN0.D XA7.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X190 AVSS XA5.XA4.MN0.G XA5.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X191 SAR_IP XB1.XA3.MN0.S XB1.XCAPB1.XCAPB4.B AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X192 XA8.XA1.XA4.MN1.D XA8.XA1.XA2.MN0.D XA8.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X193 XA0.XA4.MN0.D XA0.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X194 VREF XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X195 AVSS XB1.XA4.MN0.G XB1.XA3.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X196 AVSS CK_SAMPLE XA4.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X197 AVSS XA7.XA4.MN0.G XA7.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X198 D<0> XA8.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R23 m3_n2104_2244# XB1.XCAPB1.XCAPB4.A sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X199 VREF XA7.XA4.MN0.G XA7.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X200 AVSS XA5.XA3.MN0.G D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X201 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X202 XA8.XA1.XA1.MN0.D XA8.XA1.XA5.MN2.G XA8.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R24 XDAC1.XC0.XRES4.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X203 XA6.XA1.XA5.MN2.D EN XA6.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X204 XA4.XA1.XA4.MP1.D EN XA4.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X205 AVSS XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X206 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X207 AVSS XA0.XA12.MN0.D XA1.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X208 VREF XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R25 XDAC1.X16ab.XRES1A.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X209 XA1.XA12.MN0.G XA0.XA12.MN0.D XA1.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X210 XA6.XA4.MN0.D XA6.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X211 D<4> XA4.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X212 XA6.XA1.XA2.MN0.D XA7.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X213 AVDD EN XA4.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X214 XA5.XA9.MN1.G CK_SAMPLE XA5.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X215 XA8.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X216 XA7.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X217 XA1.XA7.MN0.D XA2.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X218 XA7.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X219 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X220 XA0.XA10.MN0.D XA0.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X221 XA1.XA7.MN0.D XA2.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X222 D<2> XA6.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X223 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X224 XA7.XA4.MN0.D XA7.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X225 XA7.XA4.MN0.D XA7.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R26 XA6.XA6.MP0.G XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X226 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X227 XA6.XA1.XA5.MP1.D EN XA6.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X228 XA6.XA9.MN0.D XA6.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X229 XA0.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R27 XDAC1.XC1.XRES1A.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X230 XA4.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X231 XA2.XA1.XA5.MN2.D XA2.XA1.XA5.MN2.G XA2.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X232 XA1.XA12.MN0.G XA1.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X233 XA1.XA11.MP0.D XA1.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X234 AVDD XA6.XA1.XA1.MN0.S XA6.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X235 XA20.XA3.MN0.D XA20.XA9.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X236 AVDD XA20.XA9.MN0.D XA20.XA3.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X237 XA2.XA4.MN0.D XA2.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X238 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X239 XA2.XA1.XA2.MN0.D XA3.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X240 SARP XB1.XA4.MN1.D SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X241 AVSS XA5.XA11.MN1.G XA5.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R28 D<8> XDAC2.XC128a<1>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X242 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X243 XA0.XA10.MN0.G XA0.XA9.MN1.G XA0.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X244 VREF XA6.XA4.MN0.G XA6.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X245 D<6> XA2.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R29 XDAC1.XC64a<0>.XRES1A.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X246 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R30 XDAC1.XC0.XRES16.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X247 XA7.XA10.MN0.D XA7.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X248 DONE XA8.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X249 XA5.XA7.MN0.D XA6.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X250 XA7.XA10.MN0.D XA7.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X251 VREF XA6.XA3.MN0.G D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X252 XA0.XA4.MN0.G EN XA0.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X253 AVSS CK_SAMPLE XA0.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X254 XA2.XA1.XA5.MN1.D XA2.XA1.XA2.MN0.D XA2.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X255 XB2.XA4.MN1.G XB2.XA1.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X256 XA8.XA6.MP0.G XA8.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X257 XA7.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X258 XA7.XA6.MP2.D D<1> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X259 SARN XB2.XA4.MN1.D SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X260 XA0.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA0.XA7.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X261 XA4.XA8.MN0.D XA4.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X262 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X263 XA5.XA12.MN0.G XA5.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X264 XA5.XA6.MP0.D XA5.XA6.MP0.G XA5.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R31 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X265 XB2.XA1.MN0.D XB2.XA1.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X266 XA6.XA9.MN1.G D<2> XA6.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X267 XA4.XA6.MP0.G XA4.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X268 AVSS XA2.XA4.MN0.G XA2.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X269 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X270 XA7.XA10.MN0.G XA7.XA9.MN1.G XA7.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X271 AVDD XA7.XA9.MN1.G XA7.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X272 AVDD XB2.XA4.MN1.D XB2.XCAPB1.XCAPB4.A AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X273 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X274 AVSS XA2.XA3.MN0.G D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X275 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X276 AVSS CK_SAMPLE XA7.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R32 XA3.XA6.MP0.G XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X277 AVDD XA7.XA6.MP0.G XA7.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R33 XA0.XA6.MP0.G XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X278 VREF XA5.XA4.MN0.D XA5.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X279 XB2.XA4.MN1.D XB2.XA4.MN1.G XB2.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X280 XA6.XA12.MN0.G XA6.XA11.MN1.G XA6.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X281 XA0.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA0.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X282 XA2.XA9.MN1.G CK_SAMPLE XA2.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X283 VREF XA5.XA4.MN0.G XA5.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X284 XA20.XA3.MN0.D SARN XA20.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X285 AVDD AVDD XA20.XA3.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R34 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X286 XA6.XA7.MN0.D XA7.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R35 XDAC1.XC64a<0>.XRES1B.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X287 VREF XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X288 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X289 AVSS XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X290 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X291 VREF XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X292 XA5.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X293 VREF XA0.XA4.MN0.D XA0.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X294 XA3.XA1.XA4.MN1.D XA3.XA1.XA2.MN0.D XA3.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X295 XA6.XA11.MP0.D XA6.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X296 XA3.XA1.XA4.MP1.D EN XA3.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X297 AVSS XA2.XA11.MN1.G XA2.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X298 XA8.XA6.MP0.D XA8.XA6.MP0.G XA8.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X299 XA5.XA4.MN0.D XA5.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R36 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X300 D<5> XA3.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X301 XA3.XA1.XA1.MN0.D XA3.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X302 VREF D<8> XA0.XA6.MP2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X303 D<5> XA3.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X304 AVDD EN XA3.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X305 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X306 AVDD XB2.XA4.MN0.G XB2.XA3.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X307 XA2.XA4.MN0.G EN XA2.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X308 XA2.XA7.MN0.D XA3.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X309 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X310 XA20.XA3.MN1.D SARN XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X311 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X312 XA20.XA3.MN6.D XA20.XA9.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X313 XB2.XA4.MN0.G CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X314 XA2.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA3.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X315 XA3.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X316 XA3.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X317 XA2.XA12.MN0.G XA2.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X318 VREF XA8.XA4.MN0.D XA8.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X319 XA5.XA10.MN0.D XA5.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R37 D<8> XDAC2.XC128a<1>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X320 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X321 XA0.XA6.MP0.G XA0.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X322 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X323 VREF XA8.XA4.MN0.G XA8.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X324 XA5.XA6.MP2.D D<3> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X325 XA4.XA1.XA5.MN2.D XA4.XA1.XA5.MN2.G XA4.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X326 VREF XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R38 XB2.XCAPB1.XCAPB4.A m3_26048_132# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X327 XB1.XA4.MN1.G XB1.XA1.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X328 XA4.XA4.MN0.D XA4.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R39 XDAC1.XC128b<2>.XRES2.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X329 XA4.XA1.XA2.MN0.D XA5.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X330 XA2.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA2.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X331 XA8.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X332 AVDD XA5.XA9.MN1.G XA5.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X333 XA3.XA8.MN0.D XA3.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X334 XA20.XA10.MN1.D XA20.XA12.MN0.D XA20.XA10.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X335 XA3.XA8.MN0.D XA3.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X336 XA6.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X337 D<4> XA4.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X338 AVDD XA20.XA12.MN0.D XA20.XA10.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X339 XA8.XA4.MN0.D XA8.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X340 AVDD XA5.XA6.MP0.G XA5.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X341 XA3.XA6.MP0.G XA3.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X342 XA3.XA6.MP0.G XA3.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X343 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R40 XDAC1.X16ab.XRES2.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X344 XA4.XA1.XA5.MN1.D XA4.XA1.XA2.MN0.D XA4.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X345 AVDD XB1.XA4.MN1.D XB1.XCAPB1.XCAPB4.A AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R41 XA5.XA6.MP0.G XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X346 XA0.XA12.MN0.D XA0.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R42 XDAC1.XC128a<1>.XRES8.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X347 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X348 VREF XA2.XA4.MN0.D XA2.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R43 D<8> XDAC2.XC128a<1>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X349 AVSS XA6.XA4.MN0.D XA6.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X350 AVSS XA4.XA4.MN0.G XA4.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X351 VREF XA2.XA3.MN0.G D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R44 XDAC1.XC1.XRES2.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R45 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X352 XA8.XA10.MN0.D XA8.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X353 AVSS XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X354 XA20.XA11.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X355 AVSS XA6.XA4.MN0.G XA6.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X356 VREF XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X357 XA20.XA11.MP0.D CK_SAMPLE AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X358 AVSS XA4.XA3.MN0.G D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X359 XA8.XA6.MP2.D D<0> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X360 XA1.XA1.XA4.MN1.D XA1.XA1.XA2.MN0.D XA1.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X361 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X362 AVSS XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X363 XA0.XA1.XA5.MN2.D EN XA0.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R46 XDAC1.XC64a<0>.XRES8.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X364 XA1.XA1.XA4.MP1.D EN XA1.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X365 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X366 D<7> XA1.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X367 XA1.XA1.XA1.MN0.D XA0.XA7.MN0.G XA1.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X368 XA0.XA4.MN0.D XA0.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X369 D<7> XA1.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X370 AVDD EN XA1.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X371 XA0.XA1.XA2.MN0.D XA0.XA7.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X372 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X373 XA4.XA9.MN1.G CK_SAMPLE XA4.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X374 XA6.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X375 XA2.XA6.MP0.G XA2.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R47 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X376 AVDD XA8.XA9.MN1.G XA8.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X377 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X378 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X379 XA6.XA4.MN0.D XA6.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X380 XA0.XA6.MP2.G D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R48 XDAC1.XC32a<0>.XRES8.B D<4> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X381 XA0.XA10.MN0.G XA0.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R49 XA2.XA3.MN0.G XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X382 AVSS XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X383 XA1.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X384 AVDD XA8.XA6.MP0.G XA8.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X385 XA0.XA1.XA5.MN1.D XA0.XA1.XA2.MN0.D XA0.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X386 XA1.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X387 XA7.XA1.XA5.MN2.D XA7.XA1.XA5.MN2.G XA7.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R50 XA3.XA3.MN0.G XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X388 XA8.XA4.MN0.G XA8.XA1.XA5.MN2.G XA8.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X389 XA7.XA1.XA5.MN2.D EN XA7.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X390 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X391 XA5.XA1.XA4.MN1.D XA5.XA1.XA2.MN0.D XA5.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X392 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X393 XA0.XA7.MN0.G XA0.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X394 AVSS XA4.XA11.MN1.G XA4.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X395 XA7.XA4.MN0.D XA7.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X396 XA7.XA4.MN0.D XA7.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X397 D<3> XA5.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X398 XA8.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X399 XA7.XA1.XA2.MN0.D XA8.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X400 XA5.XA1.XA1.MN0.D XA5.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X401 XA7.XA1.XA2.MN0.D XA8.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X402 AVSS XA0.XA4.MN0.G XA0.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X403 XA4.XA4.MN0.G EN XA4.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X404 XA6.XA10.MN0.D XA6.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X405 XA4.XA7.MN0.D XA5.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X406 D<1> XA7.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R51 XA0.XA6.MP0.G XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X407 D<1> XA7.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X408 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X409 AVSS D<8> XA0.XA6.MP2.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X410 XA4.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA5.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X411 XA3.XA11.MN1.G XA2.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X412 XA6.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X413 XA7.XA1.XA5.MN1.D XA7.XA1.XA2.MN0.D XA7.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X414 XA1.XA8.MN0.D XA1.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X415 SARN XB2.XA4.MN1.D SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X416 XA5.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X417 XA7.XA1.XA5.MP1.D EN XA7.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X418 XA1.XA8.MN0.D XA1.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X419 XA4.XA12.MN0.G XA4.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X420 XA1.XA6.MP0.G XA1.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X421 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X422 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X423 XA1.XA6.MP0.G XA1.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R52 XDAC1.XC32a<0>.XRES1A.B AVSS sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X424 AVDD XA7.XA1.XA1.MN0.S XA7.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X425 XA0.XA9.MN1.G CK_SAMPLE XA0.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X426 XA6.XA10.MN0.G XA6.XA9.MN1.G XA6.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X427 AVSS XA7.XA4.MN0.G XA7.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X428 VREF XA7.XA4.MN0.G XA7.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X429 AVSS XA20.XA2a.MN0.D XA8.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R53 XDAC1.X16ab.XRES4.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X430 AVSS CK_SAMPLE XA6.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X431 VREF XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X432 AVSS XA7.XA3.MN0.G D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X433 SARP XB1.XA4.MN1.D SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X434 VREF XA7.XA3.MN0.G D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R54 XDAC1.XC128a<1>.XRES1A.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X435 XA4.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA4.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X436 XA6.XA1.XA4.MP1.D EN XA6.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X437 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X438 XA5.XA8.MN0.D XA5.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R55 XDAC1.XC64b<1>.XRES4.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X439 AVSS XA0.XA11.MN1.G XA0.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X440 D<2> XA6.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X441 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X442 AVDD EN XA6.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X443 AVSS XA8.XA4.MN0.D XA8.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X444 XA5.XA6.MP0.G XA5.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X445 XA2.XA10.MN0.G XA2.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X446 XA7.XA9.MN1.G CK_SAMPLE XA7.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X447 XA7.XA9.MN1.G D<1> XA7.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X448 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X449 XA0.XA7.MN0.D XA0.XA7.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X450 AVSS XA8.XA3.MN0.G D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X451 AVSS XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X452 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X453 VREF XA4.XA4.MN0.D XA4.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X454 XA6.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X455 XA2.XA1.XA4.MN1.D XA2.XA1.XA2.MN0.D XA2.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R56 XDAC1.XC128b<2>.XRES4.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X456 XA0.XA12.MN0.G XA0.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X457 VREF XA4.XA3.MN0.G D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X458 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X459 D<6> XA2.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X460 XA2.XA1.XA1.MN0.D XA2.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X461 AVSS XA7.XA11.MN1.G XA7.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X462 XA7.XA12.MN0.G XA7.XA11.MN1.G XA7.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R57 XDAC1.XC32a<0>.XRES1B.B D<1> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X463 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X464 XB2.XA2.MN0.G XB2.XA2.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X465 XA8.XA6.MP0.G XA8.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X466 XA5.XA1.XA5.MN2.D EN XA5.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X467 XA7.XA7.MN0.D XA8.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X468 XA7.XA7.MN0.D XA8.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R58 D<8> XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X469 XA5.XA4.MN0.D XA5.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X470 XB2.XCAPB1.XCAPB4.B AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X471 XA2.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X472 XA5.XA1.XA2.MN0.D XA6.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X473 XA0.XA11.MN1.G XB2.XA2.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X474 XA6.XA8.MN0.D XA6.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X475 XA4.XA6.MP0.G XA4.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R59 XDAC1.XC128a<1>.XRES1B.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X476 D<3> XA5.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X477 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X478 XA7.XA12.MN0.G XA7.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X479 XB2.XCAPB1.XCAPB4.B XB2.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X480 XA7.XA11.MP0.D XA7.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X481 XA20.XA3.MN1.D SARN XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X482 XA6.XA6.MP0.G XA6.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X483 XA20.XA3.MN6.D XA20.XA3a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R60 XDAC1.XC1.XRES4.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X484 XA5.XA1.XA5.MP1.D EN XA5.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X485 XA20.XA3a.MN0.G XA20.XA3.MN6.D XA20.XA2.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X486 XA3.XA4.MN0.G XA3.XA1.XA5.MN2.G XA3.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X487 AVDD XA20.XA3.MN6.D XA20.XA3a.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X488 XA3.XA4.MN0.G EN XA3.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R61 XDAC1.XC128b<2>.XRES16.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R62 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X489 AVDD XA5.XA1.XA1.MN0.S XA5.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X490 XA0.XA6.MP0.D XA0.XA6.MP0.G XA0.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X491 XA3.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R63 XB1.XCAPB1.XCAPB4.B m3_7544_308# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X492 XA3.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA4.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X493 XA2.XA8.MN0.D XA2.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X494 VREF XA5.XA4.MN0.G XA5.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X495 XA20.XA12.MN0.G XA8.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X496 XA20.XA3.MN0.D SARN XA20.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X497 AVDD XA20.XA3a.MN0.G XA20.XA3.MN6.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X498 D<8> XA0.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R64 XB1.XCAPB1.XCAPB4.B m3_7544_3476# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X499 XA2.XA6.MP0.G XA2.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R65 XB2.XCAPB1.XCAPB4.A m3_26048_2244# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X500 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X501 AVSS XB2.XA4.MN0.G XB2.XA3.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X502 VREF XA5.XA3.MN0.G D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X503 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X504 XA5.XA11.MN1.G XA4.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X505 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X506 XA8.XA1.XA5.MN2.D EN XA8.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X507 VREF XA0.XA4.MN0.D XA0.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X508 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X509 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X510 XA8.XA4.MN0.D XA8.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X511 XA8.XA1.XA2.MN0.D XA8.XA7.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X512 XA5.XA9.MN1.G D<3> XA5.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X513 VREF XA0.XA4.MN0.G XA0.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X514 AVSS XA20.XA2a.MN0.D XA3.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X515 XA3.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA3.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X516 XA20.XA2.MN1.D SARP XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X517 D<0> XA8.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X518 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X519 XA20.XA2.MN1.D XA20.XA9.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X520 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R66 XDAC1.XC64b<1>.XRES2.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X521 AVSS XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R67 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X522 AVDD XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X523 VREF XA0.XA1.XA5.MN2.D D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R68 XA0.XA6.MP0.G XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X524 XA8.XA1.XA5.MP1.D EN XA8.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X525 XA8.XA9.MN0.D XA8.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R69 m3_16472_3476# XB2.XCAPB1.XCAPB4.B sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X526 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X527 XA0.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X528 AVSS XA3.XA4.MN0.D XA3.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X529 AVDD XA8.XA1.XA1.MN0.S XA8.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X530 XA5.XA12.MN0.G XA5.XA11.MN1.G XA5.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X531 VREF XA3.XA4.MN0.D XA3.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X532 XA20.XA12.MN0.D XA20.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X533 XA0.XA4.MN0.D XA0.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X534 XA20.XA12.MN0.D XA20.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X535 XA4.XA10.MN0.G XA4.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X536 VREF XA8.XA4.MN0.G XA8.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X537 AVSS XA3.XA3.MN0.G D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X538 XA5.XA7.MN0.D XA6.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X539 VREF XA3.XA3.MN0.G D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X540 AVDD XA20.XA9.MN0.D XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X541 AVSS XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X542 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X543 VREF XA8.XA3.MN0.G D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X544 XB1.XA2.MN0.G XB1.XA2.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X545 XA6.XA1.XA5.MN2.D XA6.XA1.XA5.MN2.G XA6.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R70 D<8> XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X546 XA20.XA4.MN0.D XA20.XA10.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X547 XA2.XA6.MP0.D XA2.XA6.MP0.G XA2.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R71 m3_n2104_1188# XB1.XCAPB1.XCAPB4.A sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X548 XA4.XA1.XA4.MN1.D XA4.XA1.XA2.MN0.D XA4.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X549 AVDD XA20.XA10.MN1.D XA20.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R72 m3_n2104_4356# XB1.XCAPB1.XCAPB4.A sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X550 XB1.XCAPB1.XCAPB4.B AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X551 XA5.XA11.MP0.D XA5.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X552 XA6.XA4.MN0.D XA6.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X553 AVSS DONE XA20.XA11.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X554 D<4> XA4.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R73 XA3.XA3.MN0.G XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X555 XA6.XA1.XA2.MN0.D XA7.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X556 XA20.XA11.MN0.D DONE XA20.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X557 XA0.XA10.MN0.D XA0.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X558 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X559 XA4.XA1.XA1.MN0.D XA4.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X560 XA8.XA9.MN1.G D<0> XA8.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X561 XA3.XA6.MP0.G XA3.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X562 XA1.XA4.MN0.G XA0.XA7.MN0.G XA1.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X563 XA3.XA6.MP0.G XA3.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X564 D<2> XA6.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X565 XA1.XA4.MN0.G EN XA1.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X566 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X567 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X568 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X569 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X570 XA0.XA6.MP2.D XA0.XA6.MP2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X571 XA1.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X572 XA20.XA3.MN6.D XA20.XA3a.MN0.G XA20.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X573 XA1.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA2.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X574 XA4.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X575 XA6.XA1.XA5.MN1.D XA6.XA1.XA2.MN0.D XA6.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X576 AVDD XA20.XA3a.MN0.G XA20.XA3.MN6.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X577 VREF XA2.XA4.MN0.D XA2.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X578 AVDD XA0.XA9.MN1.G XA0.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X579 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X580 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X581 VREF XA2.XA4.MN0.G XA2.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X582 XA8.XA12.MN0.G XA8.XA11.MN1.G XA8.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X583 AVSS XA6.XA4.MN0.G XA6.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X584 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X585 AVDD XA0.XA6.MP0.G XA0.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X586 VREF XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R74 XDAC1.XC0.XRES8.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X587 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X588 XA5.XA4.MN0.G XA5.XA1.XA5.MN2.G XA5.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X589 XA8.XA7.MN0.D XA8.XA7.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R75 D<8> XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X590 AVSS XA6.XA3.MN0.G D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X591 AVSS XA0.XA1.XA5.MN2.D D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X592 XA2.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X593 XA5.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X594 XA4.XA11.MN1.G XA3.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X595 AVSS XA20.XA2a.MN0.D XA1.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X596 XA1.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA1.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X597 XA4.XA11.MN1.G XA3.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X598 XA2.XA4.MN0.D XA2.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X599 XA0.XA1.XA4.MN1.D XA0.XA1.XA2.MN0.D XA0.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X600 XA4.XA8.MN0.D XA4.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X601 XA8.XA11.MP0.D XA8.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R76 m3_n2104_132# XB1.XCAPB1.XCAPB4.A sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X602 XA4.XA6.MP0.G XA4.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X603 XA0.XA6.MP2.G D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X604 XA0.XA1.XA1.MN0.D EN XA0.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X605 XA6.XA9.MN1.G CK_SAMPLE XA6.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X606 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X607 D<8> XA0.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X608 AVSS XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X609 VREF XA1.XA4.MN0.D XA1.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X610 AVSS XA1.XA4.MN0.D XA1.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X611 VREF XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R77 XDAC1.XC128b<2>.XRES1A.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X612 XA0.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X613 XA2.XA10.MN0.D XA2.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X614 AVSS XA1.XA3.MN0.G D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R78 m3_16472_308# XB2.XCAPB1.XCAPB4.B sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X615 XA7.XA1.XA4.MN1.D XA7.XA1.XA2.MN0.D XA7.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X616 VREF XA1.XA3.MN0.G D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X617 AVSS XA20.XA2a.MN0.D XA5.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X618 XA7.XA1.XA4.MP1.D EN XA7.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X619 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X620 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X621 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X622 AVSS XA6.XA11.MN1.G XA6.XA12.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X623 D<1> XA7.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X624 XA2.XA6.MP2.D D<6> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X625 D<1> XA7.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X626 XA7.XA1.XA1.MN0.D XA7.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X627 AVDD EN XA7.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X628 XA3.XA9.MN0.D XA3.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X629 XA6.XA4.MN0.G EN XA6.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X630 XA3.XA10.MN0.G XA3.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X631 XA6.XA7.MN0.D XA7.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X632 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R79 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X633 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X634 XA6.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA7.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X635 AVDD XA2.XA9.MN1.G XA2.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X636 XA1.XA6.MP0.G XA1.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X637 AVSS XA5.XA4.MN0.D XA5.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X638 XA7.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X639 XA1.XA6.MP0.G XA1.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X640 XA7.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X641 XA0.XA8.MN0.D XA0.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X642 XA6.XA12.MN0.G XA6.XA10.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X643 AVDD XA2.XA6.MP0.G XA2.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X644 XA8.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X645 AVSS XA5.XA3.MN0.G D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X646 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X647 XA0.XA6.MP0.G XA0.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X648 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X649 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X650 XB2.XCAPB1.XCAPB4.A XB2.XA4.MN0.G XB2.XA4.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X651 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X652 XA2.XA4.MN0.G XA2.XA1.XA5.MN2.G XA2.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X653 XA4.XA6.MP0.D XA4.XA6.MP0.G XA4.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X654 XA2.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X655 XB2.XA4.MN0.D XB2.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X656 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X657 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X658 AVSS XA8.XA4.MN0.D XA8.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X659 XA6.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA6.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X660 XA7.XA8.MN0.D XA7.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X661 XA5.XA6.MP0.G XA5.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X662 XB1.XA1.MN0.D XB1.XA1.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X663 XA7.XA8.MN0.D XA7.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R80 XDAC1.XC64a<0>.XRES4.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R81 XDAC1.XC0.XRES1A.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X664 SAR_IN XB2.XA4.MN0.G XB2.XCAPB1.XCAPB4.B AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X665 XA7.XA6.MP0.G XA7.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X666 AVSS XA8.XA4.MN0.G XA8.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X667 XA2.XA11.MN1.G XA1.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X668 XA7.XA6.MP0.G XA7.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X669 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X670 XA2.XA11.MN1.G XA1.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X671 VREF XA4.XA4.MN0.D XA4.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R82 XDAC1.X16ab.XRES16.B XA2.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X672 AVSS XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X673 SAR_IN XB2.XA3.MN0.S XB2.XCAPB1.XCAPB4.B AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X674 VREF XA6.XA4.MN0.D XA6.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X675 VREF XA4.XA4.MN0.G XA4.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R83 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X676 XB1.XA4.MN1.D XB1.XA4.MN1.G XB1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X677 AVSS XA20.XA2a.MN0.D XA2.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X678 XA8.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X679 VREF XA6.XA3.MN0.G D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X680 VREF XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R84 XDAC1.XC64b<1>.XRES16.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R85 XB1.XCAPB1.XCAPB4.B m3_7544_2420# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X681 XA8.XA4.MN0.D XA8.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X682 VREF XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R86 XA3.XA3.MN0.G XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X683 XA4.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X684 XA6.XA11.MN1.G XA5.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X685 XA5.XA1.XA4.MP1.D EN XA5.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X686 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X687 XA20.XA2.MN1.D SARP XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X688 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X689 AVSS XA2.XA4.MN0.D XA2.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X690 XA4.XA4.MN0.D XA4.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X691 XA20.XA3a.MN0.G XA20.XA9.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R87 D<8> XDAC2.XC128a<1>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X692 SARN XB2.XA4.MN1.D SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X693 D<3> XA5.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X694 AVSS XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R88 XDAC1.XC64a<0>.XRES16.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X695 AVDD EN XA5.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X696 XA1.XA9.MN0.D XA1.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X697 XA6.XA6.MP0.G XA6.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X698 AVDD XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X699 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X700 XA1.XA10.MN0.G XA1.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X701 AVSS XA2.XA3.MN0.G D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X702 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X703 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X704 XA8.XA10.MN0.D XA8.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X705 AVSS XA20.XA3.MN6.D XA20.XA2a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X706 AVDD XA20.XA3.MN6.D XA20.XA2a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X707 XA0.XA1.XA5.MN2.D EN XA0.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R89 XDAC1.XC0.XRES1B.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X708 XA5.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X709 XA8.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X710 XA0.XA4.MN0.D XA0.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R90 m3_16472_2420# XB2.XCAPB1.XCAPB4.B sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X711 XA20.XA3.MN0.D SARP XA20.XA2.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R91 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X712 XA0.XA1.XA2.MN0.D XA0.XA7.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X713 AVDD AVDD XA20.XA2.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X714 XA4.XA10.MN0.D XA4.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X715 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X716 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X717 XA0.XA6.MP2.G D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X718 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X719 XA2.XA6.MP0.G XA2.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X720 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X721 XA4.XA6.MP2.D D<4> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X722 XA8.XA10.MN0.G XA8.XA9.MN1.G XA8.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X723 XA5.XA9.MN0.D XA5.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X724 XA20.XA3.MN0.D XA20.XA9.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X725 AVDD XA20.XA9.MN0.D XA20.XA3.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X726 XA0.XA1.XA5.MP1.D EN XA0.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R92 XA4.XA6.MP0.G XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X727 XB1.XCAPB1.XCAPB4.A XB1.XA4.MN0.G XB1.XA4.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X728 AVSS CK_SAMPLE XA8.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X729 VREF XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X730 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R93 XDAC1.XC1.XRES16.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X731 XA7.XA11.MN1.G XA6.XA12.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X732 AVDD XA4.XA9.MN1.G XA4.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X733 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X734 AVDD XA0.XA1.XA1.MN0.S XA0.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R94 m3_n2104_3300# XB1.XCAPB1.XCAPB4.A sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X735 XA5.XA8.MN0.D XA5.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X736 XA3.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X737 XA8.XA1.XA4.MP1.D EN XA8.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X738 XA3.XA6.MP0.D XA3.XA6.MP0.G XA3.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X739 VREF XA0.XA4.MN0.G XA0.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X740 AVDD XA4.XA6.MP0.G XA4.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X741 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X742 XA5.XA6.MP0.G XA5.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X743 D<0> XA8.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X744 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R95 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X745 AVDD EN XA8.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X746 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X747 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X748 VREF D<8> XA0.XA6.MP2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X749 XA4.XA4.MN0.G XA4.XA1.XA5.MN2.G XA4.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X750 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X751 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X752 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X753 XB1.XA4.MN0.G CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X754 SAR_IP XB1.XA4.MN0.G XB1.XCAPB1.XCAPB4.B AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X755 XA4.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X756 XA3.XA11.MN1.G XA2.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X757 XA8.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X758 AVSS XA3.XA4.MN0.D XA3.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X759 VREF XA3.XA4.MN0.D XA3.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X760 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X761 XA0.XA9.MN1.G XA0.XA6.MP2.G XA0.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X762 AVSS XA3.XA4.MN0.G XA3.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R96 XDAC1.XC32a<0>.XRES2.B D<2> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X763 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X764 VREF XA3.XA4.MN0.G XA3.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R97 AVSS XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X765 XA20.XA10.MN0.D XA20.XA11.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X766 XA20.XA10.MN1.D XA20.XA11.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X767 XA6.XA10.MN0.G XA6.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X768 XA2.XA1.XA5.MN2.D EN XA2.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X769 AVSS XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X770 VREF XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X771 AVSS XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R98 XA3.XA3.MN0.G XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X772 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X773 XA2.XA4.MN0.D XA2.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X774 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R99 XDAC1.XC128a<1>.XRES2.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X775 XA2.XA1.XA2.MN0.D XA3.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R100 D<8> XDAC2.XC128a<1>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R101 XA0.XA6.MP0.G XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X776 XA3.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X777 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X778 XA6.XA1.XA4.MN1.D XA6.XA1.XA2.MN0.D XA6.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X779 XA3.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X780 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X781 XA0.XA12.MN0.G XA0.XA11.MN1.G XA0.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X782 D<6> XA2.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X783 AVSS XA20.XA2a.MN0.D XA4.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X784 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X785 DONE XA8.XA7.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X786 XA3.XA4.MN0.D XA3.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X787 XA3.XA4.MN0.D XA3.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X788 D<2> XA6.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R102 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X789 XA20.XA9.MN0.D XA20.XA10.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X790 XA6.XA1.XA1.MN0.D XA6.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X791 XA20.XA9.MN0.D XA20.XA10.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X792 XA0.XA7.MN0.D XA0.XA7.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X793 XA8.XA6.MP0.G XA8.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X794 XA2.XA1.XA5.MP1.D EN XA2.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X795 XA2.XA9.MN0.D XA2.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X796 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X797 SARP XB1.XA4.MN1.D SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X798 XA0.XA4.MN0.G EN XA0.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X799 AVDD XA2.XA1.XA1.MN0.S XA2.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R103 XDAC1.XC64a<0>.XRES2.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X800 AVSS XA4.XA4.MN0.D XA4.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X801 XA0.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X802 XA6.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X803 XA0.XA11.MP0.D XA0.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X804 VREF XA2.XA4.MN0.G XA2.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X805 XA3.XA10.MN0.D XA3.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R104 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X806 XA3.XA10.MN0.D XA3.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X807 AVSS XA4.XA3.MN0.G D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X808 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X809 VREF XA2.XA3.MN0.G D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R105 XDAC1.X16ab.XRES8.B XA3.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X810 XA3.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X811 XA3.XA6.MP2.D D<5> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R106 XA7.XA6.MP0.G XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X812 XA1.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X813 XA7.XA4.MN0.G XA7.XA1.XA5.MN2.G XA7.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X814 XA1.XA6.MP0.D XA1.XA6.MP0.G XA1.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X815 XA7.XA4.MN0.G EN XA7.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X816 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X817 XA7.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X818 XA2.XA9.MN1.G D<6> XA2.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X819 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X820 XA7.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA8.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X821 XA3.XA10.MN0.G XA3.XA9.MN1.G XA3.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X822 AVDD XA3.XA9.MN1.G XA3.XA10.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X823 XA6.XA8.MN0.D XA6.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X824 XA4.XA6.MP0.G XA4.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R107 D<8> XDAC2.XC128a<1>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X825 AVSS XA20.XA2a.MN0.D XA0.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X826 AVSS CK_SAMPLE XA3.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X827 XA6.XA6.MP0.G XA6.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X828 AVDD XA3.XA6.MP0.G XA3.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X829 AVSS XA1.XA4.MN0.D XA1.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X830 VREF XA1.XA4.MN0.D XA1.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X831 XA5.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X832 AVSS XA1.XA4.MN0.G XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R108 XDAC1.XC128b<2>.XRES8.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X833 XA2.XA12.MN0.G XA2.XA11.MN1.G XA2.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X834 VREF XA1.XA4.MN0.G XA1.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R109 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X835 AVSS XA0.XA4.MN0.D XA0.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X836 XA2.XA7.MN0.D XA3.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X837 AVSS XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X838 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X839 AVSS XA20.XA2a.MN0.D XA7.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X840 AVSS D<8> XA0.XA6.MP2.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X841 VREF XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X842 XA7.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA7.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X843 XA1.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R110 XB2.XCAPB1.XCAPB4.A m3_26048_1188# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X844 XA1.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X845 XA5.XA11.MN1.G XA4.XA12.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X846 XA2.XA11.MP0.D XA2.XA10.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X847 AVSS XA5.XA4.MN0.D XA5.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X848 XA1.XA4.MN0.D XA1.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X849 XA8.XA1.XA5.MN2.D XA8.XA1.XA5.MN2.G XA8.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R111 XDAC1.XC128a<1>.XRES4.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R112 XB2.XCAPB1.XCAPB4.A m3_26048_4356# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X850 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X851 XA1.XA4.MN0.D XA1.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X852 AVSS XA7.XA4.MN0.D XA7.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X853 XA8.XA4.MN0.D XA8.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X854 VREF XA7.XA4.MN0.D XA7.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X855 AVSS XA5.XA4.MN0.G XA5.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X856 XA8.XA1.XA2.MN0.D XA8.XA7.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X857 XA0.XA6.MP0.G XA0.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R113 XDAC1.XC1.XRES8.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X858 XA4.XA1.XA5.MN2.D EN XA4.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X859 AVSS XA7.XA3.MN0.G D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X860 D<0> XA8.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X861 VREF XA7.XA3.MN0.G D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X862 AVSS XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X863 XA4.XA4.MN0.D XA4.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R114 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X864 XA4.XA1.XA2.MN0.D XA5.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X865 SARP XB1.XA4.MN1.D SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X866 XA5.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X867 XA8.XA1.XA5.MN1.D XA8.XA1.XA2.MN0.D XA8.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X868 XA1.XA10.MN0.D XA1.XA10.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X869 XA1.XA10.MN0.D XA1.XA10.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X870 XA6.XA6.MP0.D XA6.XA6.MP0.G XA6.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X871 D<4> XA4.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X872 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X873 XA5.XA4.MN0.D XA5.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X874 XA0.XA11.MN1.G XB1.XA2.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X875 XA8.XA7.MN0.G XA8.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X876 XA1.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X877 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X878 XA1.XA6.MP2.D D<7> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X879 XA4.XA1.XA5.MP1.D EN XA4.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X880 XA4.XA9.MN0.D XA4.XA7.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X881 XA7.XA6.MP0.G XA7.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X882 AVSS XA8.XA4.MN0.G XA8.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X883 XA7.XA6.MP0.G XA7.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R115 XDAC1.XC32a<0>.XRES4.B D<3> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X884 XB1.XCAPB1.XCAPB4.B XB1.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X885 XA5.XA4.MN0.G EN XA5.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 SARN a_23600_51140# 0.16f
C1 XA3.XA9.MN1.G XA3.XA6.MN2.D 0.126f
C2 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES4.B 0.428f
C3 XA0.XA12.MN0.D VREF 0.39f
C4 EN a_7328_43748# 0.166f
C5 SARN XDAC2.XC1.XRES16.B 55.3f
C6 EN XA7.XA1.XA1.MN0.S 0.139f
C7 XA3.XA4.MN0.D a_7328_49028# 0.154f
C8 SARP XDAC1.XC64b<1>.XRES1A.B 3.59f
C9 XA7.XA4.MN0.G a_18560_47268# 0.157f
C10 XA5.XA1.XA5.MN2.G XA5.XA1.XA2.MN0.D 0.126f
C11 AVDD a_12368_40228# 0.464f
C12 CK_SAMPLE XA1.XA9.MN1.G 0.135f
C13 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MP1.D 0.148f
C14 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D 0.702f
C15 D<3> D<2> 6.37f
C16 AVDD a_7328_46564# 0.356f
C17 VREF D<8> 0.608f
C18 XA0.XA4.MN0.D XA1.XA3.MN0.G 0.11f
C19 AVDD a_21080_41284# 0.361f
C20 AVDD a_16040_52900# 0.387f
C21 XA1.XA3.MN0.G a_2288_46212# 0.155f
C22 XA8.XA3.MN0.G a_19928_46564# 0.156f
C23 EN a_11000_43044# 0.141f
C24 XDAC2.XC64a<0>.XRES1A.B XDAC2.XC1.XRES1B.B 0.617f
C25 XA0.XA6.MP0.G XA1.XA3.MN0.G 2.53f
C26 XA1.XA4.MN0.D SARP 0.169f
C27 AVDD XA8.XA11.MN1.G 1.04f
C28 AVDD XA8.XA7.MN0.G 5.21f
C29 XA20.XA3a.MN0.D XA5.XA1.XA2.MN0.D 0.199f
C30 XA3.XA7.MN0.D XA4.XA1.XA5.MN2.G 0.14f
C31 EN a_5960_43748# 0.166f
C32 D<3> XA7.XA6.MP0.G 0.123f
C33 D<2> XA6.XA6.MP0.G 2.21f
C34 XA7.XA4.MN0.G a_17408_47268# 0.155f
C35 AVDD a_11000_40228# 0.467f
C36 AVDD a_17408_52196# 0.37f
C37 AVDD a_2288_49732# 0.359f
C38 SARN XDAC2.XC128a<1>.XRES16.B 55.3f
C39 D<7> a_2288_50788# 0.161f
C40 AVDD a_5960_46564# 0.356f
C41 EN a_2288_42340# 0.159f
C42 D<4> XA4.XA4.MN0.G 0.26f
C43 AVDD XA2.XA1.XA2.MN0.D 0.263f
C44 SARP XDAC1.XC1.XRES16.B 55.3f
C45 XA3.XA3.MN0.G XA20.XA2a.MN0.D 0.271f
C46 AVDD a_2288_50436# 0.416f
C47 XA4.XA1.XA5.MN2.D a_11000_44452# 0.158f
C48 XA6.XA6.MP0.G XA7.XA6.MP0.G 7.36f
C49 AVDD a_17408_44452# 0.357f
C50 XA4.XA1.XA5.MN2.G XA3.XA1.XA5.MN2.D 0.108f
C51 XA0.XA6.MP0.G D<8> 5.44f
C52 AVDD XA6.XA12.MN0.G 0.709f
C53 AVDD XA8.XA1.XA5.MN2.G 4.81f
C54 AVDD a_2288_48676# 0.356f
C55 XDAC2.XC32a<0>.XRES8.B XDAC2.XC32a<0>.XRES2.B 0.44f
C56 AVDD a_17408_45508# 0.359f
C57 EN XA6.XA1.XA1.MN0.S 0.139f
C58 XA2.XA4.MN0.D a_5960_49028# 0.154f
C59 CK_SAMPLE XA0.XA9.MN1.G 0.134f
C60 AVDD a_16040_52196# 0.37f
C61 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MP1.D 0.144f
C62 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D 0.702f
C63 AVDD a_920_49732# 0.359f
C64 XB2.XCAPB1.XCAPB4.B m3_26048_2244# 0.17f
C65 EN a_920_42340# 0.159f
C66 XA2.XA3.MN0.G XA20.XA2a.MN0.D 0.26f
C67 D<8> a_920_46212# 0.155f
C68 XA7.XA3.MN0.G a_18560_46564# 0.156f
C69 XA8.XA11.MN1.G XA8.XA12.MN0.G 0.214f
C70 XB2.XCAPB1.XCAPB4.A XB2.XA4.MN0.G 0.134f
C71 AVDD a_920_50436# 0.416f
C72 SARN XDAC2.XC64b<1>.XRES16.B 55.3f
C73 XA4.XA1.XA5.MN2.D a_9848_44452# 0.153f
C74 SARN XA0.XA6.MP0.G 0.392f
C75 AVDD a_2288_47620# 0.356f
C76 XDAC1.XC64a<0>.XRES1A.B XDAC1.XC1.XRES1B.B 0.617f
C77 AVDD a_16040_44452# 0.357f
C78 AVDD a_2288_41988# 0.386f
C79 SARP XDAC1.XC128a<1>.XRES16.B 55.3f
C80 XA0.XA4.MN0.D SARP 0.391f
C81 AVDD XA7.XA11.MN1.G 1.89f
C82 AVDD a_8408_2094# 0.362f
C83 AVDD XA7.XA1.XA5.MN2.G 5.46f
C84 XA8.XA7.MN0.D a_19928_51492# 0.124f
C85 XA2.XA7.MN0.D XA3.XA1.XA5.MN2.G 0.14f
C86 AVDD a_920_48676# 0.356f
C87 AVDD a_16040_45508# 0.359f
C88 XA2.XA4.MN0.D a_4808_49028# 0.156f
C89 XA6.XA4.MN0.G a_16040_47268# 0.155f
C90 XA5.XA1.XA5.MN2.G XA4.XA1.XA2.MN0.D 0.144f
C91 SARN a_23600_49732# 0.163f
C92 D<4> D<2> 0.269f
C93 XDAC2.XC128b<2>.XRES1A.B XDAC2.XC128a<1>.XRES1B.B 0.617f
C94 AVDD XA1.XA1.XA5.MP0.D 0.159f
C95 AVDD a_17408_41284# 0.361f
C96 AVDD a_12368_52900# 0.387f
C97 XA1.XA3.MN0.G XA20.XA2a.MN0.D 0.265f
C98 D<8> a_n232_46212# 0.157f
C99 XA7.XA3.MN0.G a_17408_46564# 0.155f
C100 XA8.XA11.MN1.G XA7.XA12.MN0.G 0.391f
C101 XA20.XA4.MN0.D SARN 0.304f
C102 AVDD a_920_47620# 0.356f
C103 EN a_7328_43044# 0.141f
C104 D<0> XA8.XA4.MN0.D 0.203f
C105 XA3.XA1.XA5.MN2.G XA2.XA1.XA5.MN2.D 0.108f
C106 XA8.XA4.MN0.D XA8.XA4.MN0.G 0.708f
C107 AVDD a_920_41988# 0.386f
C108 AVDD XA5.XA12.MN0.G 0.706f
C109 XA8.XA10.MN0.D XA8.XA10.MN0.G 0.194f
C110 AVDD XB2.XCAPB1.XCAPB4.A 2.39f
C111 AVDD XA6.XA1.XA5.MN2.G 4.81f
C112 XA20.XA3a.MN0.D XA4.XA1.XA2.MN0.D 0.195f
C113 EN a_2288_43748# 0.166f
C114 SARN XDAC2.XC1.XRES2.B 6.99f
C115 SARN a_23600_48676# 0.156f
C116 D<3> XA6.XA6.MP0.G 0.121f
C117 XDAC1.XC32a<0>.XRES8.B XDAC1.XC32a<0>.XRES2.B 0.44f
C118 EN XA5.XA1.XA1.MN0.S 0.139f
C119 XA8.XA4.MN0.D a_21080_49380# 0.154f
C120 SARP XDAC1.XC64b<1>.XRES16.B 55.3f
C121 XA6.XA4.MN0.G a_14888_47268# 0.157f
C122 XA4.XA1.XA5.MN2.G XA4.XA1.XA2.MN0.D 0.126f
C123 AVDD a_7328_40228# 0.464f
C124 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D 0.702f
C125 AVDD XA20.XA3.MN0.D 0.628f
C126 AVDD a_2288_46564# 0.356f
C127 AVDD XA1.XA1.XA2.MN0.D 0.263f
C128 AVDD a_16040_41284# 0.361f
C129 AVDD a_11000_52900# 0.387f
C130 D<8> XA20.XA2a.MN0.D 0.244f
C131 XA2.XA12.MN0.G a_4808_53604# 0.1f
C132 XB2.XA4.MN1.D XB2.XA4.MN0.G 0.303f
C133 XA3.XA1.XA5.MN2.D a_8480_44452# 0.153f
C134 XDAC2.X16ab.XRES8.B XDAC2.X16ab.XRES2.B 0.44f
C135 EN a_5960_43044# 0.141f
C136 XA5.XA6.MP0.G XA7.XA6.MP0.G 0.318f
C137 AVDD XA6.XA11.MN1.G 1.04f
C138 AVDD XA5.XA1.XA5.MN2.G 5.46f
C139 XA1.XA7.MN0.D XA2.XA1.XA5.MN2.G 0.14f
C140 XA7.XA7.MN0.D a_18560_51492# 0.126f
C141 EN a_920_43748# 0.166f
C142 XA8.XA4.MN0.D a_19928_49380# 0.155f
C143 XA1.XA4.MN0.D a_3440_49028# 0.156f
C144 AVDD a_5960_40228# 0.467f
C145 AVDD a_12368_52196# 0.37f
C146 SARN XDAC2.XC128a<1>.XRES2.B 6.99f
C147 XA0.XA6.MP2.G a_920_50788# 0.161f
C148 XDAC1.XC128b<2>.XRES1A.B XDAC1.XC128a<1>.XRES1B.B 0.617f
C149 AVDD a_920_46564# 0.356f
C150 SARP a_23600_41988# 0.165f
C151 D<5> XA3.XA4.MN0.G 0.259f
C152 AVDD XA0.XA1.XA5.MP0.D 0.159f
C153 SARP XDAC1.XC1.XRES2.B 6.99f
C154 XA6.XA3.MN0.G a_16040_46564# 0.155f
C155 XA8.XA10.MN0.G XA8.XA9.MN0.D 0.106f
C156 XA7.XA11.MN1.G XA7.XA12.MN0.G 0.278f
C157 SAR_IN XB2.XCAPB1.XCAPB4.B 0.234f
C158 AVDD a_22448_50788# 0.482f
C159 XA3.XA1.XA5.MN2.D a_7328_44452# 0.158f
C160 AVDD XA20.XA3a.MN0.D 9.87f
C161 XA1.XA6.MP0.G a_2288_50084# 0.159f
C162 AVDD a_12368_44452# 0.357f
C163 XA2.XA1.XA5.MN2.G XA1.XA1.XA5.MN2.D 0.108f
C164 XA7.XA4.MN0.D XA7.XA4.MN0.G 0.707f
C165 AVDD XA4.XA12.MN0.G 0.709f
C166 XA7.XA10.MN0.D XA7.XA10.MN0.G 0.194f
C167 AVDD XB2.XA4.MN1.D 0.717f
C168 AVDD XA4.XA1.XA5.MN2.G 4.81f
C169 XA2.XA9.MN1.G XA2.XA6.MN2.D 0.126f
C170 XDAC2.XC0.XRES1A.B XDAC2.XC64b<1>.XRES1B.B 0.617f
C171 AVDD a_22448_49028# 0.488f
C172 AVDD a_12368_45508# 0.359f
C173 EN XA4.XA1.XA1.MN0.S 0.139f
C174 XA1.XA4.MN0.D a_2288_49028# 0.154f
C175 XA5.XA4.MN0.G a_13520_47268# 0.157f
C176 AVDD a_11000_52196# 0.37f
C177 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MP1.D 0.148f
C178 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D 0.702f
C179 AVDD a_22448_50084# 0.366f
C180 D<4> D<3> 5.83f
C181 XB2.XCAPB1.XCAPB4.B m3_26048_3300# 0.17f
C182 XA6.XA3.MN0.G a_14888_46564# 0.156f
C183 XA7.XA11.MN1.G XA8.XA11.MN1.G 0.271f
C184 XA8.XA10.MN0.G XA8.XA9.MN1.G 0.202f
C185 AVDD a_21080_50788# 0.361f
C186 SARN XDAC2.XC64b<1>.XRES2.B 6.99f
C187 XDAC1.X16ab.XRES8.B XDAC1.X16ab.XRES2.B 0.44f
C188 AVDD a_11000_44452# 0.357f
C189 AVDD a_22448_42340# 0.575f
C190 SARP XDAC1.XC128a<1>.XRES2.B 6.99f
C191 AVDD XA5.XA11.MN1.G 1.89f
C192 AVDD XA3.XA1.XA5.MN2.G 5.46f
C193 XA20.XA3a.MN0.D XA3.XA1.XA2.MN0.D 0.199f
C194 XA0.XA7.MN0.D XA0.XA7.MN0.G 0.14f
C195 AVDD a_21080_49028# 0.356f
C196 D<3> XA5.XA6.MP0.G 2.11f
C197 AVDD a_11000_45508# 0.359f
C198 XA7.XA4.MN0.D a_18560_49380# 0.155f
C199 XA4.XA1.XA5.MN2.G XA3.XA1.XA2.MN0.D 0.146f
C200 XA5.XA4.MN0.G a_12368_47268# 0.155f
C201 AVDD a_21080_50084# 0.361f
C202 AVDD XA8.XA3.MN0.G 2.49f
C203 XA8.XA6.MP0.G XA8.XA4.MN0.D 0.631f
C204 AVDD XA0.XA1.XA2.MN0.D 0.263f
C205 AVDD a_12368_41284# 0.361f
C206 AVDD a_7328_52900# 0.387f
C207 XA1.XA12.MN0.G a_3440_53604# 0.102f
C208 XA7.XA11.MN1.G XA6.XA12.MN0.G 0.142f
C209 XB1.XCAPB1.XCAPB4.A XB1.XA4.MN0.G 0.134f
C210 XA2.XA1.XA5.MN2.D a_5960_44452# 0.158f
C211 XA7.XA1.XA5.MN2.G XA8.XA1.XA5.MN2.G 1.58f
C212 AVDD a_22448_47972# 0.389f
C213 EN a_2288_43044# 0.141f
C214 D<1> XA7.XA4.MN0.D 0.203f
C215 XA5.XA6.MP0.G XA6.XA6.MP0.G 6.58f
C216 XA0.XA7.MN0.G XA0.XA1.XA5.MN2.D 0.108f
C217 XA6.XA4.MN0.D XA6.XA4.MN0.G 0.707f
C218 AVDD a_21080_42340# 0.361f
C219 XA6.XA10.MN0.D XA6.XA10.MN0.G 0.194f
C220 AVDD XA3.XA12.MN0.G 0.706f
C221 AVDD XB1.XCAPB1.XCAPB4.A 2.39f
C222 AVDD XA2.XA1.XA5.MN2.G 4.81f
C223 XDAC1.XC0.XRES1A.B XDAC1.XC64b<1>.XRES1B.B 0.617f
C224 SARN XDAC2.XC1.XRES8.B 27.7f
C225 EN XA3.XA1.XA1.MN0.S 0.139f
C226 XA7.XA4.MN0.D a_17408_49380# 0.154f
C227 SARP XDAC1.XC64b<1>.XRES2.B 6.99f
C228 XA3.XA1.XA5.MN2.G XA3.XA1.XA2.MN0.D 0.126f
C229 AVDD a_2288_40228# 0.464f
C230 XA0.XA7.MN0.G XA0.XA1.XA1.MP1.D 0.144f
C231 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D 0.755f
C232 XA8.XA9.MN1.G XA8.XA7.MN0.D 0.274f
C233 AVDD XA7.XA3.MN0.G 2.47f
C234 AVDD a_11000_41284# 0.361f
C235 AVDD a_5960_52900# 0.387f
C236 XA5.XA3.MN0.G a_13520_46564# 0.156f
C237 XA7.XA10.MN0.G XA7.XA9.MN0.D 0.106f
C238 XB1.XA4.MN1.D XB1.XA4.MN0.G 0.303f
C239 XA2.XA1.XA5.MN2.D a_4808_44452# 0.153f
C240 AVDD a_21080_47972# 0.356f
C241 EN a_920_43044# 0.141f
C242 XA20.XA2a.MN0.D XA8.XA1.XA1.MN0.S 0.139f
C243 XDAC2.XC64a<0>.XRES16.B XDAC2.XC64a<0>.XRES1A.B 0.454f
C244 AVDD XA4.XA11.MN1.G 1.04f
C245 AVDD XB1.XA4.MN1.D 0.717f
C246 AVDD XA0.XA7.MN0.G 5.46f
C247 XA6.XA7.MN0.D a_14888_51492# 0.124f
C248 XA0.XA4.MN0.D a_920_49028# 0.154f
C249 XA4.XA4.MN0.G a_11000_47268# 0.155f
C250 AVDD a_920_40228# 0.467f
C251 AVDD a_7328_52196# 0.37f
C252 SARN XDAC2.XC128a<1>.XRES8.B 27.7f
C253 D<6> D<2> 0.184f
C254 AVDD XA6.XA3.MN0.G 2.47f
C255 D<6> XA2.XA4.MN0.G 0.259f
C256 XA8.XA7.MN0.G XA20.XA3a.MN0.D 0.203f
C257 AVDD a_22448_43748# 0.491f
C258 SARP XDAC1.XC1.XRES8.B 27.7f
C259 XA5.XA3.MN0.G a_12368_46564# 0.155f
C260 XA7.XA10.MN0.G XA7.XA9.MN1.G 0.202f
C261 XA6.XA11.MN1.G XA6.XA12.MN0.G 0.214f
C262 SAR_IP XB1.XCAPB1.XCAPB4.B 0.234f
C263 AVDD a_17408_50788# 0.363f
C264 XA0.XA6.MP0.G a_920_50084# 0.159f
C265 AVDD a_7328_44452# 0.357f
C266 XA5.XA4.MN0.D XA5.XA4.MN0.G 0.707f
C267 AVDD XA2.XA12.MN0.G 0.709f
C268 XA5.XA10.MN0.D XA5.XA10.MN0.G 0.194f
C269 AVDD a_14960_2446# 0.406f
C270 XA20.XA3a.MN0.D XA2.XA1.XA2.MN0.D 0.195f
C271 XA1.XA9.MN1.G XA1.XA6.MN2.D 0.126f
C272 AVDD a_17408_49028# 0.356f
C273 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES8.B 0.471f
C274 AVDD a_7328_45508# 0.359f
C275 EN XA2.XA1.XA1.MN0.S 0.139f
C276 XA6.XA4.MN0.D a_16040_49380# 0.154f
C277 XA0.XA4.MN0.D a_n232_49028# 0.156f
C278 XA4.XA4.MN0.G a_9848_47268# 0.157f
C279 AVDD a_5960_52196# 0.37f
C280 XA8.XA3.MN0.G a_19928_45508# 0.104f
C281 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D 0.753f
C282 AVDD a_17408_50084# 0.358f
C283 XB2.XCAPB1.XCAPB4.B m3_26048_4356# 0.17f
C284 AVDD XA5.XA3.MN0.G 2.47f
C285 XA8.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.96f
C286 AVDD a_21080_43748# 0.357f
C287 AVDD a_16040_50788# 0.363f
C288 XA8.XA1.XA5.MN2.D a_21080_44804# 0.156f
C289 SARN XDAC2.XC64b<1>.XRES8.B 27.7f
C290 XA1.XA1.XA5.MN2.D a_3440_44452# 0.153f
C291 XA20.XA2a.MN0.D XA7.XA1.XA1.MN0.S 0.137f
C292 XA4.XA6.MP0.G XA6.XA6.MP0.G 0.321f
C293 XDAC1.XC64a<0>.XRES16.B XDAC1.XC64a<0>.XRES1A.B 0.454f
C294 AVDD a_5960_44452# 0.357f
C295 AVDD a_17408_42340# 0.361f
C296 SARP XDAC1.XC128a<1>.XRES8.B 27.7f
C297 AVDD XA3.XA11.MN1.G 1.89f
C298 AVDD a_22448_51492# 0.568f
C299 XA1.XA10.MN0.D XA1.XA10.MN0.G 0.194f
C300 XA5.XA7.MN0.D a_13520_51492# 0.126f
C301 AVDD a_16040_49028# 0.356f
C302 AVDD a_5960_45508# 0.359f
C303 XA6.XA4.MN0.D a_14888_49380# 0.155f
C304 XA8.XA7.MN0.G XA8.XA3.MN0.G 0.106f
C305 XA3.XA1.XA5.MN2.G XA2.XA1.XA2.MN0.D 0.144f
C306 XA7.XA9.MN1.G XA7.XA7.MN0.D 0.274f
C307 AVDD a_16040_50084# 0.358f
C308 XDAC2.XC128b<2>.XRES16.B XDAC2.XC128b<2>.XRES1A.B 0.454f
C309 AVDD XA4.XA3.MN0.G 2.47f
C310 XA7.XA6.MP0.G XA7.XA4.MN0.D 0.76f
C311 XA7.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.885f
C312 AVDD a_7328_41284# 0.361f
C313 AVDD a_2288_52900# 0.387f
C314 XA4.XA3.MN0.G a_11000_46564# 0.155f
C315 XA6.XA11.MN1.G XA5.XA12.MN0.G 0.391f
C316 XA6.XA10.MN0.G XA6.XA9.MN0.D 0.106f
C317 XA8.XA1.XA5.MN2.D a_19928_44804# 0.153f
C318 XA1.XA1.XA5.MN2.D a_2288_44452# 0.158f
C319 XA5.XA1.XA5.MN2.G XA6.XA1.XA5.MN2.G 1.58f
C320 AVDD a_17408_47972# 0.356f
C321 D<2> XA6.XA4.MN0.D 0.203f
C322 D<0> VREF 1.29f
C323 XA4.XA4.MN0.D XA4.XA4.MN0.G 0.707f
C324 VREF XA8.XA4.MN0.G 0.258f
C325 AVDD a_16040_42340# 0.361f
C326 AVDD XA1.XA12.MN0.G 0.706f
C327 XA4.XA10.MN0.D XA4.XA10.MN0.G 0.194f
C328 AVDD a_21080_51492# 0.387f
C329 SARN XDAC2.XC1.XRES4.B 13.9f
C330 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES8.B 0.471f
C331 EN XA1.XA1.XA1.MN0.S 0.139f
C332 SARP XDAC1.XC64b<1>.XRES8.B 27.7f
C333 XA2.XA1.XA5.MN2.G XA2.XA1.XA2.MN0.D 0.126f
C334 XA3.XA4.MN0.G a_8480_47268# 0.157f
C335 AVDD a_22448_40580# 0.483f
C336 XA7.XA3.MN0.G a_18560_45508# 0.106f
C337 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D 0.755f
C338 D<5> D<4> 0.348f
C339 AVDD XA3.XA3.MN0.G 2.47f
C340 XA6.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.963f
C341 AVDD a_5960_41284# 0.361f
C342 AVDD a_920_52900# 0.387f
C343 XA4.XA3.MN0.G a_9848_46564# 0.156f
C344 XA0.XA12.MN0.G a_n232_53604# 0.1f
C345 XA6.XA10.MN0.G XA6.XA9.MN1.G 0.202f
C346 XB2.XA4.MN1.D XB2.XCAPB1.XCAPB4.A 0.233f
C347 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES8.B 0.471f
C348 AVDD a_16040_47972# 0.356f
C349 XA20.XA2a.MN0.D XA6.XA1.XA1.MN0.S 0.137f
C350 EN a_21080_43396# 0.162f
C351 XA20.XA3.MN0.D XA20.XA3a.MN0.D 0.176f
C352 VREF XA7.XA4.MN0.G 0.263f
C353 AVDD XA2.XA11.MN1.G 1.04f
C354 XA0.XA10.MN0.D XA0.XA10.MN0.G 0.194f
C355 XA20.XA3a.MN0.D XA1.XA1.XA2.MN0.D 0.199f
C356 XA8.XA4.MN0.G XA8.XA1.XA2.MN0.D 0.206f
C357 D<4> XA4.XA6.MP0.G 2.1f
C358 XA8.XA1.XA5.MN2.G XA7.XA3.MN0.G 0.106f
C359 XA5.XA4.MN0.D a_13520_49380# 0.155f
C360 AVDD a_22448_43044# 0.419f
C361 XA3.XA4.MN0.G a_7328_47268# 0.155f
C362 AVDD a_21080_40580# 0.381f
C363 AVDD a_2288_52196# 0.37f
C364 XA0.XA4.MN0.G EN 0.227f
C365 SARN XDAC2.XC128a<1>.XRES4.B 13.9f
C366 XDAC1.XC128b<2>.XRES16.B XDAC1.XC128b<2>.XRES1A.B 0.454f
C367 AVDD XA2.XA3.MN0.G 2.47f
C368 D<7> XA1.XA4.MN0.G 0.259f
C369 XA5.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.885f
C370 AVDD a_17408_43748# 0.357f
C371 SARP XDAC1.XC1.XRES4.B 13.9f
C372 XA5.XA11.MN1.G XA5.XA12.MN0.G 0.278f
C373 XB2.XA4.MN1.D XB2.XA4.MN0.D 0.139f
C374 AVDD a_12368_50788# 0.363f
C375 XA7.XA1.XA5.MN2.D a_18560_44804# 0.153f
C376 XA0.XA1.XA5.MN2.D a_920_44452# 0.158f
C377 XA4.XA6.MP0.G XA5.XA6.MP0.G 6.62f
C378 AVDD a_2288_44452# 0.357f
C379 XA3.XA4.MN0.D XA3.XA4.MN0.G 0.728f
C380 VREF XA6.XA4.MN0.G 0.263f
C381 AVDD XA0.XA12.MN0.G 0.709f
C382 XA3.XA10.MN0.D XA3.XA10.MN0.G 0.194f
C383 XDAC2.XC0.XRES16.B XDAC2.XC0.XRES1A.B 0.454f
C384 AVDD a_12368_49028# 0.356f
C385 AVDD a_2288_45508# 0.359f
C386 EN XA0.XA1.XA1.MN0.S 0.17f
C387 XA5.XA4.MN0.D a_12368_49380# 0.154f
C388 AVDD a_21080_43044# 0.381f
C389 AVDD a_920_52196# 0.37f
C390 D<8> XA0.XA1.XA5.MN2.D 0.753f
C391 XA6.XA9.MN1.G XA6.XA7.MN0.D 0.274f
C392 AVDD a_12368_50084# 0.358f
C393 AVDD XA1.XA3.MN0.G 2.47f
C394 XA4.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.963f
C395 AVDD a_16040_43748# 0.357f
C396 AVDD XA20.XA9.MN0.D 4.02f
C397 XA3.XA3.MN0.G a_8480_46564# 0.156f
C398 XA5.XA11.MN1.G XA6.XA11.MN1.G 0.271f
C399 XA5.XA10.MN0.G XA5.XA9.MN0.D 0.106f
C400 AVDD a_11000_50788# 0.363f
C401 XA7.XA1.XA5.MN2.D a_17408_44804# 0.156f
C402 XA0.XA1.XA5.MN2.D a_n232_44452# 0.153f
C403 SARN XDAC2.XC64b<1>.XRES4.B 13.9f
C404 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES8.B 0.471f
C405 XA20.XA2a.MN0.D XA5.XA1.XA1.MN0.S 0.137f
C406 D<1> VREF 1.3f
C407 AVDD a_920_44452# 0.357f
C408 VREF XA5.XA4.MN0.G 0.263f
C409 AVDD a_12368_42340# 0.361f
C410 SARP XDAC1.XC128a<1>.XRES4.B 13.9f
C411 AVDD XA0.XA12.MN0.D 1.89f
C412 AVDD a_8408_2446# 0.406f
C413 AVDD a_17408_51492# 0.387f
C414 XA4.XA7.MN0.D a_9848_51492# 0.124f
C415 AVDD a_11000_49028# 0.356f
C416 AVDD a_920_45508# 0.359f
C417 XA7.XA1.XA5.MN2.G XA6.XA3.MN0.G 0.106f
C418 XA2.XA1.XA5.MN2.G XA1.XA1.XA2.MN0.D 0.146f
C419 XA2.XA4.MN0.G a_5960_47268# 0.155f
C420 XA20.XA10.MN1.D XA20.XA9.MN0.D 2.14f
C421 SARN a_23600_52196# 0.156f
C422 AVDD a_11000_50084# 0.358f
C423 D<6> D<4> 0.568f
C424 XB2.XCAPB1.XCAPB4.A m3_16472_308# 0.106f
C425 AVDD D<8> 2.47f
C426 XA20.XA3a.MN0.G a_22448_49732# 0.159f
C427 XA8.XA6.MP0.G VREF 0.5f
C428 XA3.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.885f
C429 XA6.XA6.MP0.G XA6.XA4.MN0.D 0.76f
C430 XA20.XA3.MN6.D XA20.XA2a.MN0.D 0.431f
C431 AVDD a_2288_41284# 0.361f
C432 AVDD XA8.XA10.MN0.D 0.728f
C433 XA3.XA3.MN0.G a_7328_46564# 0.155f
C434 XA5.XA11.MN1.G XA4.XA12.MN0.G 0.142f
C435 AVDD XA1.XA10.MN0.D 0.727f
C436 XA5.XA10.MN0.G XA5.XA9.MN1.G 0.202f
C437 SAR_IN XB2.XA4.MN0.G 0.115f
C438 XA3.XA1.XA5.MN2.G XA4.XA1.XA5.MN2.G 1.58f
C439 AVDD a_12368_47972# 0.356f
C440 EN a_17408_43396# 0.162f
C441 D<3> XA5.XA4.MN0.D 0.203f
C442 XA2.XA4.MN0.D XA2.XA4.MN0.G 0.728f
C443 XA20.XA3a.MN0.G a_23600_47620# 0.154f
C444 VREF XA4.XA4.MN0.G 0.263f
C445 AVDD a_11000_42340# 0.361f
C446 XA8.XA10.MN0.D a_19928_52900# 0.128f
C447 XA2.XA10.MN0.D XA2.XA10.MN0.G 0.194f
C448 AVDD XB2.XA4.MN1.G 0.433f
C449 AVDD a_16040_51492# 0.387f
C450 XA20.XA3a.MN0.D XA0.XA1.XA2.MN0.D 0.195f
C451 XA0.XA9.MN1.G XA0.XA6.MN2.D 0.126f
C452 XDAC1.XC0.XRES16.B XDAC1.XC0.XRES1A.B 0.454f
C453 SARN XDAC2.XC1.XRES1B.B 3.59f
C454 D<3> XA2.XA6.MP0.G 0.191f
C455 D<1> XA0.XA6.MP0.G 0.173f
C456 XA4.XA4.MN0.D a_11000_49380# 0.154f
C457 SARP XDAC1.XC64b<1>.XRES4.B 13.9f
C458 XA0.XA7.MN0.G XA1.XA1.XA2.MN0.D 0.126f
C459 XA2.XA4.MN0.G a_4808_47268# 0.157f
C460 AVDD a_17408_40580# 0.381f
C461 AVDD SARN 0.139f
C462 XA6.XA3.MN0.G a_14888_45508# 0.104f
C463 XA0.XA11.MN1.G CK_SAMPLE_BSSW 4.96f
C464 SARP a_23600_44452# 0.154f
C465 XA2.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.963f
C466 XA20.XA3a.MN0.G XA20.XA2a.MN0.D 0.222f
C467 AVDD a_920_41284# 0.361f
C468 AVDD XA7.XA10.MN0.D 0.727f
C469 AVDD XA0.XA10.MN0.D 0.728f
C470 XA6.XA1.XA5.MN2.D a_16040_44804# 0.156f
C471 AVDD a_11000_47972# 0.356f
C472 XA20.XA2a.MN0.D XA4.XA1.XA1.MN0.S 0.137f
C473 EN a_16040_43396# 0.162f
C474 XDAC2.XC64a<0>.XRES2.B XDAC2.XC64a<0>.XRES16.B 0.457f
C475 AVDD SARP 0.16f
C476 XA20.XA3a.MN0.G a_22448_47620# 0.181f
C477 VREF XA3.XA4.MN0.G 0.263f
C478 AVDD a_22448_53956# 0.405f
C479 XA20.XA10.MN1.D SARN 0.869f
C480 XA7.XA4.MN0.G XA7.XA1.XA2.MN0.D 0.206f
C481 XA3.XA7.MN0.D a_8480_51492# 0.126f
C482 XA6.XA1.XA5.MN2.G XA5.XA3.MN0.G 0.106f
C483 XA4.XA4.MN0.D a_9848_49380# 0.155f
C484 AVDD a_17408_43044# 0.381f
C485 XA8.XA4.MN0.G a_21080_47620# 0.155f
C486 AVDD a_16040_40580# 0.381f
C487 XA5.XA9.MN1.G XA5.XA7.MN0.D 0.274f
C488 SARN XDAC2.XC128a<1>.XRES1B.B 3.59f
C489 XB1.XCAPB1.XCAPB4.B m3_n2104_132# 0.17f
C490 AVDD a_22448_46916# 0.363f
C491 XA0.XA6.MP2.G XA0.XA4.MN0.G 0.259f
C492 XA0.XA7.MN0.G XA20.XA3a.MN0.D 0.885f
C493 AVDD a_12368_43748# 0.357f
C494 XA20.XA10.MN1.D SARP 0.423f
C495 SARP XDAC1.XC1.XRES1B.B 3.59f
C496 AVDD XA6.XA10.MN0.D 0.728f
C497 XA2.XA3.MN0.G a_5960_46564# 0.155f
C498 XA8.XA4.MN0.G XA8.XA1.XA5.MN2.D 0.135f
C499 XA4.XA10.MN0.G XA4.XA9.MN0.D 0.106f
C500 XA4.XA11.MN1.G XA4.XA12.MN0.G 0.214f
C501 AVDD a_7328_50788# 0.363f
C502 XA6.XA1.XA5.MN2.D a_14888_44804# 0.153f
C503 D<2> VREF 1.3f
C504 XA1.XA4.MN0.D XA1.XA4.MN0.G 0.728f
C505 VREF XA2.XA4.MN0.G 0.263f
C506 AVDD a_21080_53956# 0.461f
C507 XA7.XA10.MN0.D a_18560_52900# 0.13f
C508 AVDD XB2.XA1.MN0.D 0.514f
C509 AVDD a_7328_49028# 0.356f
C510 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES4.B 0.428f
C511 AVDD a_22448_45860# 0.403f
C512 SARP a_23600_41284# 0.16f
C513 AVDD a_16040_43044# 0.381f
C514 XA1.XA4.MN0.G a_3440_47268# 0.157f
C515 XA8.XA4.MN0.G a_19928_47620# 0.154f
C516 AVDD XA8.XA9.MN1.G 0.926f
C517 XA5.XA3.MN0.G a_13520_45508# 0.106f
C518 AVDD a_7328_50084# 0.358f
C519 D<6> D<5> 0.832f
C520 AVDD a_21080_46916# 0.359f
C521 XA7.XA6.MP0.G VREF 0.568f
C522 AVDD a_11000_43748# 0.357f
C523 AVDD XA8.XA1.XA1.MP2.D 0.127f
C524 AVDD XA5.XA10.MN0.D 0.727f
C525 XA2.XA3.MN0.G a_4808_46564# 0.156f
C526 XA4.XA10.MN0.G XA4.XA9.MN1.G 0.202f
C527 AVDD a_22448_53252# 0.388f
C528 XB1.XA4.MN1.D XB1.XA4.MN0.D 0.139f
C529 SAR_IP XB1.XA4.MN0.G 0.115f
C530 AVDD a_5960_50788# 0.363f
C531 SARN XDAC2.XC64b<1>.XRES1B.B 3.59f
C532 XA20.XA2a.MN0.D XA3.XA1.XA1.MN0.S 0.137f
C533 XDAC1.XC64a<0>.XRES2.B XDAC1.XC64a<0>.XRES16.B 0.457f
C534 AVDD a_22448_44804# 0.366f
C535 VREF XA1.XA4.MN0.G 0.263f
C536 AVDD a_7328_42340# 0.361f
C537 SARP XDAC1.XC128a<1>.XRES1B.B 3.59f
C538 AVDD a_12368_51492# 0.387f
C539 AVDD a_5960_49028# 0.356f
C540 D<3> XA1.XA6.MP0.G 0.11f
C541 D<5> XA3.XA6.MP0.G 0.537f
C542 AVDD a_21080_45860# 0.356f
C543 XA3.XA4.MN0.D a_8480_49380# 0.155f
C544 XA5.XA1.XA5.MN2.G XA4.XA3.MN0.G 0.106f
C545 XA0.XA7.MN0.G XA0.XA1.XA2.MN0.D 0.144f
C546 XA1.XA4.MN0.G a_2288_47268# 0.155f
C547 AVDD a_5960_50084# 0.358f
C548 XB2.XCAPB1.XCAPB4.A m3_16472_1364# 0.106f
C549 XDAC2.XC128b<2>.XRES2.B XDAC2.XC128b<2>.XRES16.B 0.457f
C550 XA5.XA6.MP0.G XA5.XA4.MN0.D 0.76f
C551 XA8.XA6.MP0.G a_21080_49732# 0.101f
C552 AVDD XA8.XA1.XA1.MN0.S 1.05f
C553 AVDD XA4.XA10.MN0.D 0.728f
C554 XA7.XA4.MN0.G XA7.XA1.XA5.MN2.D 0.135f
C555 XA4.XA11.MN1.G XA3.XA12.MN0.G 0.391f
C556 AVDD a_21080_53252# 0.364f
C557 XB1.XA4.MN1.D XB1.XCAPB1.XCAPB4.A 0.233f
C558 XA5.XA1.XA5.MN2.D a_13520_44804# 0.153f
C559 XA0.XA7.MN0.G XA2.XA1.XA5.MN2.G 1.58f
C560 AVDD a_7328_47972# 0.356f
C561 EN a_12368_43396# 0.162f
C562 XA3.XA6.MP0.G XA4.XA6.MP0.G 4.3f
C563 D<4> XA4.XA4.MN0.D 0.203f
C564 AVDD a_21080_44804# 0.356f
C565 VREF XA0.XA4.MN0.G 0.263f
C566 AVDD a_5960_42340# 0.361f
C567 AVDD XB1.XA1.MN0.D 0.514f
C568 AVDD a_11000_51492# 0.387f
C569 SARN XDAC2.XC64a<0>.XRES1A.B 3.59f
C570 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES4.B 0.428f
C571 XA3.XA4.MN0.D a_7328_49380# 0.154f
C572 SARP XDAC1.XC64b<1>.XRES1B.B 3.59f
C573 XA7.XA4.MN0.G a_18560_47620# 0.154f
C574 AVDD a_12368_40580# 0.381f
C575 AVDD XA7.XA9.MN1.G 0.93f
C576 XA4.XA9.MN1.G XA4.XA7.MN0.D 0.274f
C577 AVDD XA7.XA1.XA1.MP2.D 0.127f
C578 AVDD XA3.XA10.MN0.D 0.727f
C579 XA1.XA3.MN0.G a_3440_46564# 0.156f
C580 XA3.XA10.MN0.G XA3.XA9.MN0.D 0.106f
C581 XA5.XA1.XA5.MN2.D a_12368_44804# 0.156f
C582 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES4.B 0.428f
C583 AVDD a_5960_47972# 0.356f
C584 XA20.XA2a.MN0.D XA2.XA1.XA1.MN0.S 0.137f
C585 EN a_11000_43396# 0.162f
C586 D<3> VREF 1.3f
C587 D<4> XA3.XA4.MN0.D 3.22f
C588 XA0.XA4.MN0.D XA0.XA4.MN0.G 0.728f
C589 XA20.XA3a.MN0.D XA3.XA3.MN0.G 0.223f
C590 AVDD a_17408_53956# 0.464f
C591 AVDD XB1.XA4.MN1.G 0.433f
C592 XA6.XA4.MN0.G XA6.XA1.XA2.MN0.D 0.206f
C593 XA7.XA7.MN0.D XA7.XA8.MN0.D 0.124f
C594 XA2.XA7.MN0.D a_4808_51492# 0.124f
C595 CK_SAMPLE VREF 1.93f
C596 XA4.XA1.XA5.MN2.G XA3.XA3.MN0.G 0.225f
C597 AVDD a_12368_43044# 0.381f
C598 XA0.XA4.MN0.G a_920_47268# 0.155f
C599 XA7.XA4.MN0.G a_17408_47620# 0.155f
C600 AVDD a_11000_40580# 0.381f
C601 SARN XDAC2.XC128b<2>.XRES1A.B 3.59f
C602 D<7> D<5> 0.146f
C603 XB1.XCAPB1.XCAPB4.B m3_n2104_1188# 0.17f
C604 XDAC1.XC128b<2>.XRES2.B XDAC1.XC128b<2>.XRES16.B 0.457f
C605 AVDD a_17408_46916# 0.359f
C606 XA6.XA6.MP0.G VREF 0.568f
C607 AVDD a_7328_43748# 0.357f
C608 AVDD XA7.XA1.XA1.MN0.S 1.03f
C609 SARP XDAC1.XC64a<0>.XRES1A.B 3.59f
C610 AVDD XA2.XA10.MN0.D 0.728f
C611 XA1.XA3.MN0.G a_2288_46564# 0.155f
C612 XA6.XA4.MN0.G XA6.XA1.XA5.MN2.D 0.135f
C613 XA3.XA11.MN1.G XA3.XA12.MN0.G 0.278f
C614 XA3.XA10.MN0.G XA3.XA9.MN1.G 0.202f
C615 AVDD a_2288_50788# 0.363f
C616 XA20.XA9.MN0.D XA20.XA3.MN0.D 0.35f
C617 D<4> XA2.XA4.MN0.D 0.192f
C618 XA20.XA3a.MN0.D XA2.XA3.MN0.G 0.221f
C619 XA6.XA10.MN0.D a_14888_52900# 0.128f
C620 AVDD a_16040_53956# 0.461f
C621 AVDD a_14960_2798# 0.465f
C622 XDAC2.XC0.XRES2.B XDAC2.XC0.XRES16.B 0.457f
C623 AVDD a_2288_49028# 0.356f
C624 D<3> XA0.XA6.MP0.G 0.102f
C625 AVDD a_17408_45860# 0.356f
C626 XA2.XA4.MN0.D a_5960_49380# 0.154f
C627 XA3.XA1.XA5.MN2.G XA3.XA3.MN0.G 0.229f
C628 AVDD a_11000_43044# 0.381f
C629 XA0.XA4.MN0.G a_n232_47268# 0.157f
C630 AVDD XA6.XA9.MN1.G 0.93f
C631 XA4.XA3.MN0.G a_9848_45508# 0.104f
C632 AVDD a_2288_50084# 0.358f
C633 AVDD a_16040_46916# 0.359f
C634 AVDD a_5960_43748# 0.357f
C635 AVDD XA6.XA1.XA1.MP2.D 0.127f
C636 XA3.XA11.MN1.G XA4.XA11.MN1.G 0.271f
C637 AVDD a_17408_53252# 0.361f
C638 AVDD a_920_50788# 0.363f
C639 XA4.XA1.XA5.MN2.D a_11000_44804# 0.156f
C640 SARN XDAC2.XC0.XRES1A.B 3.59f
C641 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES4.B 0.428f
C642 XA20.XA2a.MN0.D XA1.XA1.XA1.MN0.S 0.137f
C643 AVDD a_17408_44804# 0.356f
C644 AVDD a_2288_42340# 0.361f
C645 SARP XDAC1.XC128b<2>.XRES1A.B 3.59f
C646 XA20.XA3a.MN0.D XA1.XA3.MN0.G 0.219f
C647 AVDD a_7328_51492# 0.387f
C648 SARN XB2.XCAPB1.XCAPB4.A 1.53f
C649 XA6.XA7.MN0.D XA6.XA8.MN0.D 0.124f
C650 XA1.XA7.MN0.D a_3440_51492# 0.126f
C651 AVDD a_920_49028# 0.356f
C652 AVDD a_16040_45860# 0.356f
C653 XA2.XA4.MN0.D a_4808_49380# 0.155f
C654 XA3.XA1.XA5.MN2.G XA2.XA3.MN0.G 0.12f
C655 XA6.XA4.MN0.G a_16040_47620# 0.155f
C656 XA8.XA7.MN0.G XA8.XA1.XA1.MN0.S 0.305f
C657 XA3.XA9.MN1.G XA3.XA7.MN0.D 0.274f
C658 AVDD a_920_50084# 0.358f
C659 SARN XA20.XA3.MN0.D 0.422f
C660 XB2.XCAPB1.XCAPB4.A m3_16472_2420# 0.106f
C661 XA4.XA6.MP0.G XA4.XA4.MN0.D 0.76f
C662 AVDD XA6.XA1.XA1.MN0.S 1.04f
C663 D<8> a_920_46564# 0.155f
C664 XA5.XA4.MN0.G XA5.XA1.XA5.MN2.D 0.135f
C665 XA3.XA11.MN1.G XA2.XA12.MN0.G 0.142f
C666 AVDD a_16040_53252# 0.364f
C667 XA2.XA10.MN0.G XA2.XA9.MN0.D 0.106f
C668 XA4.XA1.XA5.MN2.D a_9848_44804# 0.153f
C669 AVDD a_2288_47972# 0.356f
C670 EN a_7328_43396# 0.162f
C671 D<5> XA3.XA4.MN0.D 7.46f
C672 D<4> VREF 1.3f
C673 AVDD a_16040_44804# 0.356f
C674 AVDD a_920_42340# 0.361f
C675 XA20.XA3.MN0.D SARP 0.511f
C676 XA20.XA3a.MN0.D D<8> 0.207f
C677 XA5.XA10.MN0.D a_13520_52900# 0.13f
C678 AVDD a_5960_51492# 0.387f
C679 XDAC1.XC0.XRES2.B XDAC1.XC0.XRES16.B 0.457f
C680 SARN XDAC2.XC64a<0>.XRES16.B 55.3f
C681 SARN a_23600_49028# 0.156f
C682 XA2.XA1.XA5.MN2.G XA2.XA3.MN0.G 0.326f
C683 SARP XDAC1.XC0.XRES1A.B 3.59f
C684 XA6.XA4.MN0.G a_14888_47620# 0.154f
C685 AVDD a_7328_40580# 0.381f
C686 AVDD XA5.XA9.MN1.G 0.93f
C687 XA3.XA3.MN0.G a_8480_45508# 0.109f
C688 XA0.XA6.MP2.G D<5> 0.185f
C689 D<7> D<6> 1.33f
C690 XA5.XA6.MP0.G VREF 0.568f
C691 AVDD XA5.XA1.XA1.MP2.D 0.127f
C692 D<8> a_n232_46564# 0.156f
C693 XA2.XA10.MN0.G XA2.XA9.MN1.G 0.202f
C694 XB2.XA4.MN1.G XB2.XA4.MN1.D 0.129f
C695 AVDD XA8.XA6.MP2.D 0.163f
C696 AVDD a_920_47972# 0.356f
C697 XA20.XA2a.MN0.D XA0.XA1.XA1.MN0.S 0.137f
C698 EN a_5960_43396# 0.162f
C699 D<5> XA2.XA4.MN0.D 3.83f
C700 XDAC2.XC64a<0>.XRES8.B XDAC2.XC64a<0>.XRES2.B 0.44f
C701 AVDD a_12368_53956# 0.464f
C702 SARN XB2.XA4.MN1.D 0.285f
C703 XA5.XA4.MN0.G XA5.XA1.XA2.MN0.D 0.206f
C704 XA5.XA7.MN0.D XA5.XA8.MN0.D 0.124f
C705 D<6> XA2.XA6.MP0.G 0.468f
C706 XA1.XA4.MN0.D a_3440_49380# 0.155f
C707 XA2.XA1.XA5.MN2.G XA1.XA3.MN0.G 0.222f
C708 AVDD a_7328_43044# 0.381f
C709 AVDD a_5960_40580# 0.381f
C710 AVDD XA20.XA3.MN1.D 0.439f
C711 SARN XDAC2.XC128b<2>.XRES16.B 55.3f
C712 XB1.XCAPB1.XCAPB4.B m3_n2104_2244# 0.17f
C713 AVDD a_12368_46916# 0.359f
C714 EN a_21080_42692# 0.159f
C715 AVDD a_2288_43748# 0.357f
C716 AVDD XA5.XA1.XA1.MN0.S 1.03f
C717 SARP XDAC1.XC64a<0>.XRES16.B 55.3f
C718 XA4.XA4.MN0.G XA4.XA1.XA5.MN2.D 0.135f
C719 XA2.XA11.MN1.G XA2.XA12.MN0.G 0.214f
C720 AVDD a_14960_n18# 0.445f
C721 SAR_IN XB2.XA4.MN1.D 0.682f
C722 XA3.XA1.XA5.MN2.D a_8480_44804# 0.153f
C723 XA2.XA6.MP0.G XA3.XA6.MP0.G 1.9f
C724 D<5> XA1.XA4.MN0.D 0.267f
C725 AVDD XA20.XA1.MN0.D 0.478f
C726 DONE CK_SAMPLE 0.155f
C727 AVDD a_11000_53956# 0.461f
C728 AVDD a_22448_49380# 0.368f
C729 XDAC2.XC128a<1>.XRES1A.B XDAC2.XC32a<0>.XRES1B.B 0.617f
C730 AVDD a_12368_45860# 0.356f
C731 XA1.XA4.MN0.D a_2288_49380# 0.154f
C732 XA0.XA7.MN0.G XA1.XA3.MN0.G 0.229f
C733 AVDD a_5960_43044# 0.381f
C734 XA20.XA3.MN6.D a_23600_45508# 0.154f
C735 XA5.XA4.MN0.G a_13520_47620# 0.154f
C736 AVDD XA4.XA9.MN1.G 0.93f
C737 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.S 0.301f
C738 XA2.XA9.MN1.G XA2.XA7.MN0.D 0.274f
C739 CK_SAMPLE a_19928_50436# 0.161f
C740 AVDD XA20.XA3.MN6.D 5.96f
C741 AVDD a_11000_46916# 0.359f
C742 AVDD a_920_43748# 0.357f
C743 XA20.XA10.MN1.D XA20.XA1.MN0.D 0.112f
C744 AVDD XA4.XA1.XA1.MP2.D 0.127f
C745 XA1.XA10.MN0.G XA1.XA9.MN0.D 0.106f
C746 XA8.XA10.MN0.G a_19928_52548# 0.128f
C747 AVDD a_12368_53252# 0.361f
C748 AVDD D<0> 2.26f
C749 XA3.XA1.XA5.MN2.D a_7328_44804# 0.156f
C750 SARN XDAC2.XC0.XRES16.B 55.3f
C751 AVDD XA8.XA4.MN0.G 2.39f
C752 D<5> VREF 1.3f
C753 XDAC1.XC64a<0>.XRES8.B XDAC1.XC64a<0>.XRES2.B 0.44f
C754 AVDD a_12368_44804# 0.356f
C755 AVDD XA8.XA1.XA4.MP0.D 0.147f
C756 SARP XDAC1.XC128b<2>.XRES16.B 55.3f
C757 XA20.XA3.MN6.D a_22448_44452# 0.16f
C758 AVDD a_8408_2798# 0.464f
C759 AVDD a_2288_51492# 0.387f
C760 XA20.XA2a.MN0.D XA20.XA2.MN1.D 0.103f
C761 XA4.XA7.MN0.D XA4.XA8.MN0.D 0.124f
C762 XA0.XA7.MN0.D a_n232_51492# 0.124f
C763 AVDD a_21080_49380# 0.356f
C764 XA20.XA10.MN1.D XA20.XA3.MN6.D 0.196f
C765 AVDD a_11000_45860# 0.356f
C766 XA0.XA7.MN0.G D<8> 0.12f
C767 XA20.XA3.MN6.D a_22448_45508# 0.168f
C768 XA5.XA4.MN0.G a_12368_47620# 0.155f
C769 CK_SAMPLE a_18560_50436# 0.161f
C770 AVDD XA20.XA3a.MN0.G 5.77f
C771 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128b<2>.XRES2.B 0.44f
C772 XB2.XCAPB1.XCAPB4.A m3_16472_3476# 0.106f
C773 XA3.XA6.MP0.G XA3.XA4.MN0.D 4.49f
C774 XA4.XA6.MP0.G VREF 0.568f
C775 SARP XB1.XCAPB1.XCAPB4.A 1.54f
C776 AVDD XA4.XA1.XA1.MN0.S 1.04f
C777 XA3.XA4.MN0.G XA3.XA1.XA5.MN2.D 0.135f
C778 XA2.XA11.MN1.G XA1.XA12.MN0.G 0.391f
C779 AVDD a_11000_53252# 0.364f
C780 XA1.XA10.MN0.G XA1.XA9.MN1.G 0.202f
C781 AVDD XA7.XA4.MN0.G 2.36f
C782 EN a_2288_43396# 0.162f
C783 D<6> XA2.XA4.MN0.D 7.43f
C784 D<5> XA0.XA4.MN0.D 0.455f
C785 AVDD a_11000_44804# 0.356f
C786 XA4.XA10.MN0.D a_9848_52900# 0.128f
C787 AVDD a_14960_3150# 0.485f
C788 AVDD a_920_51492# 0.387f
C789 SARN XB1.XA4.MN1.D 0.141f
C790 XA20.XA10.MN1.D XA20.XA3a.MN0.G 0.15f
C791 SARP a_23600_43748# 0.155f
C792 SARN XDAC2.XC64a<0>.XRES2.B 6.99f
C793 XDAC1.XC128a<1>.XRES1A.B XDAC1.XC32a<0>.XRES1B.B 0.617f
C794 SARP XDAC1.XC0.XRES16.B 55.3f
C795 AVDD a_2288_40580# 0.381f
C796 AVDD XA3.XA9.MN1.G 0.93f
C797 XA2.XA3.MN0.G a_4808_45508# 0.107f
C798 AVDD XA8.XA6.MP0.D 0.157f
C799 EN a_17408_42692# 0.159f
C800 SARP XB1.XA4.MN1.D 0.228f
C801 AVDD XA3.XA1.XA1.MP2.D 0.127f
C802 XA2.XA3.MN0.G XA3.XA3.MN0.G 1.48f
C803 XA7.XA10.MN0.G a_18560_52548# 0.13f
C804 AVDD XA7.XA6.MP2.D 0.172f
C805 XA2.XA1.XA5.MN2.D a_5960_44804# 0.156f
C806 XDAC2.XC64b<1>.XRES1A.B XDAC2.X16ab.XRES1B.B 0.617f
C807 AVDD XA6.XA4.MN0.G 2.36f
C808 EN a_920_43396# 0.162f
C809 D<6> XA1.XA4.MN0.D 6.17f
C810 AVDD a_7328_53956# 0.464f
C811 XA1.XA10.MN0.D a_3440_52900# 0.13f
C812 XA4.XA4.MN0.G XA4.XA1.XA2.MN0.D 0.206f
C813 XA3.XA7.MN0.D XA3.XA8.MN0.D 0.124f
C814 SARN a_23600_51492# 0.157f
C815 XA0.XA4.MN0.D a_920_49380# 0.154f
C816 AVDD a_2288_43044# 0.381f
C817 XA4.XA4.MN0.G a_11000_47620# 0.155f
C818 AVDD a_920_40580# 0.381f
C819 XA8.XA3.MN0.G a_21080_45860# 0.155f
C820 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S 0.327f
C821 XA1.XA9.MN1.G XA1.XA7.MN0.D 0.274f
C822 SARN XDAC2.XC128b<2>.XRES2.B 6.99f
C823 XB1.XCAPB1.XCAPB4.B m3_n2104_3300# 0.17f
C824 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128b<2>.XRES2.B 0.44f
C825 AVDD a_7328_46916# 0.359f
C826 EN a_16040_42692# 0.159f
C827 XA6.XA6.MP0.G a_16040_49732# 0.101f
C828 AVDD XA3.XA1.XA1.MN0.S 1.03f
C829 SARP XDAC1.XC64a<0>.XRES2.B 6.99f
C830 XA1.XA3.MN0.G XA3.XA3.MN0.G 0.171f
C831 XA2.XA4.MN0.G XA2.XA1.XA5.MN2.D 0.135f
C832 XA0.XA12.MN0.D XA1.XA12.MN0.G 0.278f
C833 XA0.XA10.MN0.G XA0.XA9.MN0.D 0.106f
C834 AVDD D<1> 2.31f
C835 XA2.XA1.XA5.MN2.D a_4808_44804# 0.153f
C836 AVDD XA5.XA4.MN0.G 2.36f
C837 D<6> VREF 1.3f
C838 AVDD XA7.XA1.XA4.MP0.D 0.152f
C839 AVDD a_5960_53956# 0.461f
C840 XA3.XA10.MN0.D a_8480_52900# 0.13f
C841 AVDD XB2.XA2.MN0.G 0.788f
C842 AVDD XA7.XA8.MN0.D 0.227f
C843 XA8.XA7.MN0.D a_21080_51844# 0.133f
C844 XDAC2.XC0.XRES8.B XDAC2.XC0.XRES2.B 0.44f
C845 AVDD a_17408_49380# 0.356f
C846 XA8.XA7.MN0.G XA20.XA3.MN6.D 0.256f
C847 AVDD a_7328_45860# 0.356f
C848 VREF XA8.XA4.MN0.D 0.588f
C849 XA0.XA4.MN0.D a_n232_49380# 0.155f
C850 AVDD a_920_43044# 0.381f
C851 XA4.XA4.MN0.G a_9848_47620# 0.154f
C852 AVDD XA2.XA9.MN1.G 0.93f
C853 XA1.XA3.MN0.G a_3440_45508# 0.109f
C854 XA8.XA3.MN0.G a_19928_45860# 0.162f
C855 CK_SAMPLE a_14888_50436# 0.161f
C856 AVDD XA8.XA6.MP0.G 1.65f
C857 XA0.XA6.MP2.G D<7> 2.22f
C858 XA8.XA7.MN0.G D<0> 0.6f
C859 AVDD a_5960_46916# 0.359f
C860 XA8.XA7.MN0.G XA8.XA4.MN0.G 0.158f
C861 XA3.XA6.MP0.G VREF 0.568f
C862 XA20.XA9.MN0.D a_22448_43044# 0.139f
C863 AVDD XA2.XA1.XA1.MP2.D 0.127f
C864 D<8> XA3.XA3.MN0.G 0.216f
C865 XA1.XA3.MN0.G XA2.XA3.MN0.G 3.47f
C866 XA0.XA12.MN0.D XA2.XA11.MN1.G 0.271f
C867 XA0.XA10.MN0.G XA0.XA9.MN1.G 0.202f
C868 AVDD a_7328_53252# 0.361f
C869 AVDD a_8408_n18# 0.444f
C870 SAR_IP XB1.XA4.MN1.D 0.679f
C871 AVDD XA6.XA6.MP2.D 0.172f
C872 SARN XDAC2.XC0.XRES2.B 6.99f
C873 XDAC1.XC64b<1>.XRES1A.B XDAC1.X16ab.XRES1B.B 0.617f
C874 AVDD XA4.XA4.MN0.G 2.36f
C875 D<6> XA0.XA4.MN0.D 0.293f
C876 AVDD a_7328_44804# 0.356f
C877 AVDD XA6.XA1.XA4.MP0.D 0.152f
C878 SARP XDAC1.XC128b<2>.XRES2.B 6.99f
C879 XA20.XA12.MN0.D CK_SAMPLE 0.155f
C880 AVDD a_14960_3502# 0.468f
C881 AVDD XA6.XA8.MN0.D 0.227f
C882 XA2.XA7.MN0.D XA2.XA8.MN0.D 0.124f
C883 XA8.XA7.MN0.D a_19928_51844# 0.159f
C884 AVDD a_16040_49380# 0.356f
C885 D<7> XA1.XA6.MP0.G 0.537f
C886 AVDD a_5960_45860# 0.356f
C887 VREF XA7.XA4.MN0.D 0.593f
C888 CK_SAMPLE a_13520_50436# 0.161f
C889 XB2.XCAPB1.XCAPB4.A m3_16472_4532# 0.106f
C890 XA2.XA6.MP0.G XA2.XA4.MN0.D 4.49f
C891 XA8.XA1.XA5.MN2.G XA8.XA4.MN0.G 0.168f
C892 XDAC2.XC1.XRES16.B XDAC2.XC1.XRES1A.B 0.454f
C893 AVDD XA2.XA1.XA1.MN0.S 1.04f
C894 VREF EN 0.911f
C895 XA1.XA4.MN0.G XA1.XA1.XA5.MN2.D 0.135f
C896 AVDD a_5960_53252# 0.364f
C897 XA0.XA12.MN0.D XA0.XA12.MN0.G 0.142f
C898 AVDD a_14960_334# 0.486f
C899 XA1.XA1.XA5.MN2.D a_3440_44804# 0.153f
C900 XA8.XA1.XA5.MN2.D a_21080_45156# 0.155f
C901 AVDD XA3.XA4.MN0.G 2.36f
C902 D<7> XA1.XA4.MN0.D 6.79f
C903 XA1.XA6.MP0.G XA2.XA6.MP0.G 2.62f
C904 AVDD a_5960_44804# 0.356f
C905 AVDD XA5.XA8.MN0.D 0.227f
C906 XDAC1.XC0.XRES8.B XDAC1.XC0.XRES2.B 0.44f
C907 SARN XDAC2.XC64a<0>.XRES8.B 27.7f
C908 VREF XA6.XA4.MN0.D 0.593f
C909 SARP XDAC1.XC0.XRES2.B 6.99f
C910 XA3.XA4.MN0.G a_8480_47620# 0.154f
C911 AVDD a_22448_40932# 0.57f
C912 AVDD XA1.XA9.MN1.G 0.93f
C913 XA7.XA3.MN0.G a_18560_45860# 0.162f
C914 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.S 0.301f
C915 XA0.XA9.MN1.G XA0.XA7.MN0.D 0.274f
C916 AVDD XA7.XA6.MP0.D 0.144f
C917 EN a_12368_42692# 0.159f
C918 XA8.XA1.XA5.MN2.G XA7.XA4.MN0.G 0.158f
C919 XA20.XA3.MN1.D XA20.XA3.MN0.D 0.547f
C920 AVDD XA1.XA1.XA1.MP2.D 0.127f
C921 D<8> XA1.XA3.MN0.G 3.29f
C922 XA6.XA10.MN0.G a_14888_52548# 0.128f
C923 XB1.XA4.MN1.G XB1.XA4.MN1.D 0.129f
C924 AVDD D<2> 2.31f
C925 XA1.XA1.XA5.MN2.D a_2288_44804# 0.156f
C926 XA8.XA1.XA5.MN2.D a_19928_45156# 0.153f
C927 AVDD XA2.XA4.MN0.G 2.36f
C928 D<7> VREF 1.3f
C929 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES8.B 0.471f
C930 AVDD a_2288_53956# 0.464f
C931 AVDD a_14960_3854# 0.447f
C932 XA0.XA10.MN0.D a_n232_52900# 0.128f
C933 AVDD XA4.XA8.MN0.D 0.227f
C934 XA3.XA4.MN0.G XA3.XA1.XA2.MN0.D 0.206f
C935 XA1.XA7.MN0.D XA1.XA8.MN0.D 0.124f
C936 XA7.XA7.MN0.D a_18560_51844# 0.159f
C937 VREF XA5.XA4.MN0.D 0.593f
C938 XA2.XA4.MN0.D XA3.XA4.MN0.D 0.935f
C939 AVDD a_22448_43396# 0.438f
C940 XA3.XA4.MN0.G a_7328_47620# 0.155f
C941 AVDD a_21080_40932# 0.358f
C942 XA7.XA3.MN0.G a_17408_45860# 0.155f
C943 AVDD XA7.XA6.MP0.G 6.09f
C944 SARN XDAC2.XC128b<2>.XRES8.B 27.7f
C945 XB1.XCAPB1.XCAPB4.B m3_n2104_4356# 0.17f
C946 AVDD a_2288_46916# 0.359f
C947 EN a_11000_42692# 0.159f
C948 XA7.XA1.XA5.MN2.G XA7.XA4.MN0.G 0.169f
C949 SARN XA1.XA3.MN0.G 0.137f
C950 XA20.XA3.MN6.D XA20.XA3.MN0.D 0.338f
C951 XA2.XA6.MP0.G VREF 0.568f
C952 XDAC1.XC1.XRES16.B XDAC1.XC1.XRES1A.B 0.454f
C953 AVDD XA1.XA1.XA1.MN0.S 1.03f
C954 SARP XDAC1.XC64a<0>.XRES8.B 27.7f
C955 XA0.XA4.MN0.G XA0.XA1.XA5.MN2.D 0.135f
C956 XA20.XA9.MN0.D SARN 0.652f
C957 AVDD XA1.XA4.MN0.G 2.36f
C958 D<7> XA0.XA4.MN0.D 2.87f
C959 AVDD XA5.XA1.XA4.MP0.D 0.152f
C960 AVDD a_920_53956# 0.461f
C961 XA2.XA10.MN0.D a_4808_52900# 0.128f
C962 AVDD XA3.XA8.MN0.D 0.227f
C963 XA7.XA7.MN0.D a_17408_51844# 0.133f
C964 AVDD a_12368_49380# 0.356f
C965 XDAC2.XC128a<1>.XRES16.B XDAC2.XC128a<1>.XRES1A.B 0.454f
C966 AVDD a_2288_45860# 0.356f
C967 VREF XA4.XA4.MN0.D 0.593f
C968 XA20.XA9.MN0.D SARP 0.405f
C969 AVDD a_21080_43396# 0.36f
C970 AVDD XA0.XA9.MN1.G 0.93f
C971 D<8> a_n232_45508# 0.107f
C972 CK_SAMPLE a_9848_50436# 0.161f
C973 AVDD XA6.XA6.MP0.D 0.144f
C974 XA8.XA1.XA5.MN2.G D<1> 0.704f
C975 AVDD a_920_46916# 0.359f
C976 XA7.XA1.XA5.MN2.G XA6.XA4.MN0.G 0.158f
C977 SARN D<8> 0.327f
C978 XA20.XA3a.MN0.G XA20.XA3.MN0.D 0.357f
C979 AVDD XA0.XA1.XA1.MP2.D 0.127f
C980 XA5.XA10.MN0.G a_13520_52548# 0.13f
C981 AVDD a_2288_53252# 0.361f
C982 AVDD XA5.XA6.MP2.D 0.172f
C983 SARN XDAC2.XC0.XRES8.B 27.7f
C984 XA0.XA1.XA5.MN2.D a_920_44804# 0.156f
C985 XA7.XA1.XA5.MN2.D a_18560_45156# 0.153f
C986 AVDD XA0.XA4.MN0.G 2.36f
C987 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES8.B 0.471f
C988 AVDD a_2288_44804# 0.356f
C989 XA20.XA3.MN6.D XA20.XA3a.MN0.D 0.449f
C990 XA8.XA4.MN0.D a_21080_48676# 0.154f
C991 AVDD XA4.XA1.XA4.MP0.D 0.152f
C992 SARP XDAC1.XC128b<2>.XRES8.B 27.7f
C993 AVDD XA2.XA8.MN0.D 0.227f
C994 D<8> SARP 0.2f
C995 XA0.XA7.MN0.D XA0.XA8.MN0.D 0.124f
C996 AVDD a_11000_49380# 0.356f
C997 AVDD a_920_45860# 0.356f
C998 VREF XA3.XA4.MN0.D 0.615f
C999 XA1.XA4.MN0.D XA2.XA4.MN0.D 1.55f
C1000 XA2.XA4.MN0.G a_5960_47620# 0.155f
C1001 XA6.XA3.MN0.G a_16040_45860# 0.155f
C1002 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S 0.327f
C1003 CK_SAMPLE a_8480_50436# 0.161f
C1004 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES8.B 0.471f
C1005 XA6.XA1.XA5.MN2.G XA6.XA4.MN0.G 0.168f
C1006 XA1.XA6.MP0.G XA1.XA4.MN0.D 4.65f
C1007 AVDD XA0.XA1.XA1.MN0.S 1.04f
C1008 AVDD a_920_53252# 0.364f
C1009 AVDD D<3> 2.31f
C1010 XA0.XA1.XA5.MN2.D a_n232_44804# 0.153f
C1011 XA7.XA1.XA5.MN2.D a_17408_45156# 0.155f
C1012 XA20.XA2a.MN0.D EN 0.897f
C1013 XA0.XA6.MP2.G VREF 1.3f
C1014 AVDD a_920_44804# 0.356f
C1015 SARN SARP 6.27f
C1016 XA20.XA3a.MN0.G XA20.XA3a.MN0.D 0.515f
C1017 XA8.XA4.MN0.D a_19928_48676# 0.158f
C1018 AVDD CK_SAMPLE 5.8f
C1019 AVDD a_8408_3150# 0.487f
C1020 AVDD XA1.XA8.MN0.D 0.227f
C1021 SARN SAR_IN 1.01f
C1022 XA6.XA7.MN0.D a_16040_51844# 0.133f
C1023 SARN XDAC2.XC64a<0>.XRES4.B 13.9f
C1024 D<0> a_21080_50788# 0.161f
C1025 XDAC1.XC128a<1>.XRES16.B XDAC1.XC128a<1>.XRES1A.B 0.454f
C1026 VREF XA2.XA4.MN0.D 0.615f
C1027 SARP XDAC1.XC0.XRES8.B 27.7f
C1028 XA7.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C1029 XA2.XA4.MN0.G a_4808_47620# 0.154f
C1030 AVDD a_17408_40932# 0.358f
C1031 AVDD a_22448_52548# 0.573f
C1032 XA6.XA3.MN0.G a_14888_45860# 0.162f
C1033 XB2.XA4.MN0.G CK_SAMPLE_BSSW 0.148f
C1034 AVDD XA6.XA6.MP0.G 5.96f
C1035 EN a_7328_42692# 0.159f
C1036 XA6.XA1.XA5.MN2.G XA5.XA4.MN0.G 0.158f
C1037 XA0.XA6.MP0.G XA3.XA4.MN0.D 0.869f
C1038 XA20.XA3a.MN0.G a_22448_50084# 0.156f
C1039 XA1.XA6.MP0.G VREF 0.568f
C1040 SARP SAR_IN 0.606f
C1041 AVDD a_8408_334# 0.487f
C1042 XB2.XA1.MN0.D XB2.XA4.MN1.G 0.208f
C1043 AVDD XA4.XA6.MP2.D 0.172f
C1044 XDAC2.XC64b<1>.XRES16.B XDAC2.XC64b<1>.XRES1A.B 0.454f
C1045 AVDD a_22448_48324# 0.416f
C1046 XA0.XA6.MP2.G XA0.XA4.MN0.D 9.98f
C1047 D<0> XA8.XA3.MN0.G 0.534f
C1048 XA8.XA4.MN0.G XA8.XA3.MN0.G 0.554f
C1049 AVDD XB1.XA2.MN0.G 0.788f
C1050 AVDD XA0.XA8.MN0.D 0.227f
C1051 XA2.XA4.MN0.G XA2.XA1.XA2.MN0.D 0.206f
C1052 XA6.XA7.MN0.D a_14888_51844# 0.159f
C1053 XA0.XA6.MP2.G XA0.XA6.MP0.G 0.468f
C1054 VREF XA1.XA4.MN0.D 0.615f
C1055 AVDD a_17408_43396# 0.361f
C1056 XA6.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C1057 AVDD a_16040_40932# 0.358f
C1058 AVDD a_21080_52548# 0.405f
C1059 XB2.XA4.MN0.G a_14960_686# 0.119f
C1060 XB1.XA4.MN0.G CK_SAMPLE_BSSW 0.148f
C1061 XA8.XA1.XA5.MN2.D EN 0.122f
C1062 SARN XDAC2.XC128b<2>.XRES4.B 13.9f
C1063 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES8.B 0.471f
C1064 AVDD a_22448_47268# 0.404f
C1065 EN a_5960_42692# 0.159f
C1066 XA5.XA1.XA5.MN2.G XA5.XA4.MN0.G 0.169f
C1067 XA0.XA6.MP0.G XA2.XA4.MN0.D 0.412f
C1068 AVDD a_22448_41636# 0.569f
C1069 SARP XDAC1.XC64a<0>.XRES4.B 13.9f
C1070 AVDD XA8.XA11.MP0.D 0.19f
C1071 AVDD CK_SAMPLE_BSSW 14.7f
C1072 XA6.XA1.XA5.MN2.D a_16040_45156# 0.155f
C1073 AVDD a_21080_48324# 0.359f
C1074 XA0.XA6.MP0.G XA1.XA6.MP0.G 6.08f
C1075 AVDD XA20.XA2.MN1.D 0.461f
C1076 XA7.XA4.MN0.D a_18560_48676# 0.158f
C1077 AVDD XA3.XA1.XA4.MP0.D 0.152f
C1078 AVDD a_22448_54308# 0.364f
C1079 SARN SAR_IP 0.683f
C1080 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES8.B 0.471f
C1081 AVDD a_7328_49380# 0.356f
C1082 XA8.XA1.XA5.MN2.G XA7.XA6.MP0.G 0.185f
C1083 AVDD a_22448_46212# 0.368f
C1084 XA0.XA4.MN0.D XA1.XA4.MN0.D 4.7f
C1085 AVDD a_16040_43396# 0.361f
C1086 XA1.XA4.MN0.G a_3440_47620# 0.154f
C1087 XA5.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C1088 XA8.XA4.MN0.G a_21080_47972# 0.155f
C1089 XA5.XA3.MN0.G a_13520_45860# 0.162f
C1090 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.S 0.301f
C1091 XB2.XA4.MN0.G a_13808_686# 0.113f
C1092 AVDD XA5.XA6.MP0.D 0.144f
C1093 CK_SAMPLE a_4808_50436# 0.161f
C1094 XA7.XA1.XA5.MN2.D EN 0.121f
C1095 XA7.XA1.XA5.MN2.G D<2> 0.627f
C1096 XB1.XCAPB1.XCAPB4.A m3_7544_308# 0.106f
C1097 AVDD a_21080_47268# 0.356f
C1098 XA0.XA6.MP0.G XA1.XA4.MN0.D 0.294f
C1099 XA5.XA1.XA5.MN2.G XA4.XA4.MN0.G 0.158f
C1100 SARP SAR_IP 1.01f
C1101 AVDD a_21080_41636# 0.404f
C1102 AVDD XA7.XA11.MP0.D 0.176f
C1103 XA4.XA10.MN0.G a_9848_52548# 0.128f
C1104 AVDD a_14960_686# 0.37f
C1105 AVDD D<4> 2.31f
C1106 SARN XDAC2.XC0.XRES4.B 13.9f
C1107 XA6.XA1.XA5.MN2.D a_14888_45156# 0.153f
C1108 XDAC1.XC64b<1>.XRES16.B XDAC1.XC64b<1>.XRES1A.B 0.454f
C1109 XA7.XA4.MN0.D a_17408_48676# 0.154f
C1110 AVDD XA2.XA1.XA4.MP0.D 0.152f
C1111 SARP XDAC1.XC128b<2>.XRES4.B 13.9f
C1112 XA7.XA4.MN0.G XA7.XA3.MN0.G 0.554f
C1113 AVDD a_21080_54308# 0.447f
C1114 AVDD a_8408_3502# 0.467f
C1115 AVDD a_22448_51844# 0.568f
C1116 XA5.XA7.MN0.D a_13520_51844# 0.159f
C1117 AVDD a_5960_49380# 0.356f
C1118 XA7.XA1.XA5.MN2.G XA7.XA6.MP0.G 0.149f
C1119 AVDD a_21080_46212# 0.356f
C1120 XA0.XA4.MN0.D VREF 0.615f
C1121 XA1.XA4.MN0.G a_2288_47620# 0.155f
C1122 XA4.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C1123 XA8.XA4.MN0.G a_19928_47972# 0.153f
C1124 XA5.XA3.MN0.G a_12368_45860# 0.155f
C1125 AVDD XA5.XA6.MP0.G 5.95f
C1126 CK_SAMPLE a_3440_50436# 0.161f
C1127 XA6.XA1.XA5.MN2.D EN 0.122f
C1128 XA4.XA1.XA5.MN2.G XA4.XA4.MN0.G 0.168f
C1129 XA4.XA6.MP0.G a_11000_49732# 0.101f
C1130 XA0.XA6.MP0.G VREF 0.568f
C1131 XDAC2.XC1.XRES2.B XDAC2.XC1.XRES16.B 0.457f
C1132 AVDD XA6.XA11.MP0.D 0.19f
C1133 AVDD a_22448_45156# 0.405f
C1134 AVDD a_21080_51844# 0.385f
C1135 XA5.XA7.MN0.D a_12368_51844# 0.133f
C1136 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES8.B 0.471f
C1137 SARN XDAC2.XC64a<0>.XRES1B.B 3.59f
C1138 SARP XDAC1.XC0.XRES4.B 13.9f
C1139 XA3.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C1140 AVDD a_12368_40932# 0.358f
C1141 AVDD a_17408_52548# 0.405f
C1142 AVDD XA4.XA6.MP0.D 0.144f
C1143 XA5.XA1.XA5.MN2.D EN 0.121f
C1144 XA8.XA1.XA5.MN2.D a_21080_44100# 0.126f
C1145 EN a_2288_42692# 0.159f
C1146 XA8.XA6.MP0.G a_21080_50084# 0.159f
C1147 XA0.XA6.MP0.G XA0.XA4.MN0.D 4.81f
C1148 XA4.XA1.XA5.MN2.G XA3.XA4.MN0.G 0.158f
C1149 XA3.XA10.MN0.G a_8480_52548# 0.13f
C1150 AVDD XA5.XA11.MP0.D 0.176f
C1151 AVDD XA3.XA6.MP2.D 0.172f
C1152 XA5.XA1.XA5.MN2.D a_13520_45156# 0.153f
C1153 AVDD a_17408_48324# 0.359f
C1154 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES4.B 0.428f
C1155 AVDD a_21080_45156# 0.356f
C1156 XA6.XA4.MN0.D a_16040_48676# 0.154f
C1157 D<1> XA7.XA3.MN0.G 0.572f
C1158 XA6.XA4.MN0.G XA6.XA3.MN0.G 0.554f
C1159 AVDD a_8408_3854# 0.448f
C1160 XA1.XA4.MN0.G XA1.XA1.XA2.MN0.D 0.206f
C1161 AVDD a_12368_43396# 0.361f
C1162 XA0.XA4.MN0.G a_920_47620# 0.155f
C1163 XA2.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C1164 XA7.XA4.MN0.G a_18560_47972# 0.153f
C1165 AVDD a_11000_40932# 0.358f
C1166 AVDD a_16040_52548# 0.405f
C1167 XA4.XA3.MN0.G a_11000_45860# 0.155f
C1168 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S 0.327f
C1169 XA0.XA11.MN1.G a_12368_1742# 0.156f
C1170 SARN XDAC2.XC128b<2>.XRES1B.B 3.59f
C1171 XA4.XA1.XA5.MN2.D EN 0.122f
C1172 AVDD a_17408_47268# 0.356f
C1173 EN a_920_42692# 0.159f
C1174 XA3.XA1.XA5.MN2.G XA3.XA4.MN0.G 0.169f
C1175 XDAC1.XC1.XRES2.B XDAC1.XC1.XRES16.B 0.457f
C1176 AVDD a_17408_41636# 0.404f
C1177 SARP XDAC1.XC64a<0>.XRES1B.B 3.59f
C1178 AVDD XA4.XA11.MP0.D 0.19f
C1179 AVDD D<5> 2.23f
C1180 XA5.XA1.XA5.MN2.D a_12368_45156# 0.155f
C1181 AVDD a_16040_48324# 0.359f
C1182 XA6.XA4.MN0.D a_14888_48676# 0.158f
C1183 AVDD XA1.XA1.XA4.MP0.D 0.152f
C1184 AVDD a_17408_54308# 0.448f
C1185 XA4.XA7.MN0.D a_11000_51844# 0.133f
C1186 AVDD a_2288_49380# 0.356f
C1187 D<1> a_17408_50788# 0.161f
C1188 XDAC2.XC128a<1>.XRES2.B XDAC2.XC128a<1>.XRES16.B 0.457f
C1189 AVDD a_17408_46212# 0.356f
C1190 AVDD a_11000_43396# 0.361f
C1191 XA1.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C1192 XA0.XA4.MN0.G a_n232_47620# 0.154f
C1193 XA7.XA4.MN0.G a_17408_47972# 0.155f
C1194 XA4.XA3.MN0.G a_9848_45860# 0.162f
C1195 XA0.XA11.MN1.G a_11000_1742# 0.155f
C1196 XB1.XA4.MN0.G a_9560_686# 0.114f
C1197 XB2.XA4.MN1.D a_12368_334# 0.157f
C1198 CK_SAMPLE a_n232_50436# 0.161f
C1199 AVDD XA4.XA6.MP0.G 5.98f
C1200 XA3.XA1.XA5.MN2.D EN 0.121f
C1201 XA6.XA1.XA5.MN2.G D<3> 0.704f
C1202 XB1.XCAPB1.XCAPB4.A m3_7544_1364# 0.106f
C1203 AVDD a_16040_47268# 0.356f
C1204 XA3.XA1.XA5.MN2.G XA2.XA4.MN0.G 0.158f
C1205 AVDD a_16040_41636# 0.404f
C1206 AVDD XA3.XA11.MP0.D 0.176f
C1207 AVDD XA2.XA6.MP2.D 0.172f
C1208 SARN XDAC2.XC0.XRES1B.B 3.62f
C1209 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES4.B 0.428f
C1210 AVDD XA0.XA1.XA4.MP0.D 0.152f
C1211 SARP XDAC1.XC128b<2>.XRES1B.B 3.59f
C1212 XA5.XA4.MN0.G XA5.XA3.MN0.G 0.554f
C1213 AVDD a_16040_54308# 0.447f
C1214 AVDD a_22448_39876# 0.438f
C1215 AVDD a_17408_51844# 0.387f
C1216 XA4.XA7.MN0.D a_9848_51844# 0.159f
C1217 DONE VREF 0.108f
C1218 AVDD a_920_49380# 0.356f
C1219 SARN XDAC2.XC32a<0>.XRES1A.B 3.59f
C1220 AVDD a_16040_46212# 0.356f
C1221 XA0.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C1222 XA8.XA7.MN0.G a_19928_41636# 0.128f
C1223 XB1.XA4.MN0.G a_8408_686# 0.118f
C1224 XA20.XA2a.MN0.D XA8.XA1.XA2.MN0.D 0.225f
C1225 XA2.XA1.XA5.MN2.D EN 0.122f
C1226 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES4.B 0.428f
C1227 XA2.XA1.XA5.MN2.G XA2.XA4.MN0.G 0.168f
C1228 AVDD XA2.XA11.MP0.D 0.19f
C1229 AVDD a_8408_686# 0.37f
C1230 XB1.XA4.MN1.G XB1.XA1.MN0.D 0.208f
C1231 XA4.XA1.XA5.MN2.D a_11000_45156# 0.155f
C1232 XA20.XA9.MN0.D XA20.XA3.MN6.D 0.343f
C1233 AVDD a_17408_45156# 0.356f
C1234 XA5.XA4.MN0.D a_13520_48676# 0.158f
C1235 VREF XA8.XA1.XA5.MN2.D 0.336f
C1236 AVDD a_21080_39876# 0.44f
C1237 AVDD a_16040_51844# 0.387f
C1238 SARN a_23600_49380# 0.157f
C1239 XDAC1.XC128a<1>.XRES2.B XDAC1.XC128a<1>.XRES16.B 0.457f
C1240 SARP XDAC1.XC0.XRES1B.B 3.6f
C1241 XA6.XA4.MN0.G a_16040_47972# 0.155f
C1242 AVDD a_7328_40932# 0.358f
C1243 AVDD a_12368_52548# 0.405f
C1244 XA3.XA3.MN0.G a_8480_45860# 0.162f
C1245 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MN0.S 0.301f
C1246 XB2.XA4.MN0.G a_13808_1038# 0.158f
C1247 AVDD XA3.XA6.MP0.D 0.144f
C1248 XA7.XA1.XA5.MN2.D a_17408_44100# 0.124f
C1249 XA1.XA1.XA5.MN2.D EN 0.121f
C1250 SARN XA20.XA3.MN1.D 0.143f
C1251 XA2.XA1.XA5.MN2.G XA1.XA4.MN0.G 0.158f
C1252 XA2.XA10.MN0.G a_4808_52548# 0.128f
C1253 AVDD XA1.XA11.MP0.D 0.176f
C1254 AVDD a_14960_1038# 0.489f
C1255 AVDD D<6> 2.23f
C1256 XA4.XA1.XA5.MN2.D a_9848_45156# 0.153f
C1257 XA20.XA9.MN0.D XA20.XA3a.MN0.G 0.519f
C1258 XDAC2.XC64b<1>.XRES2.B XDAC2.XC64b<1>.XRES16.B 0.457f
C1259 AVDD a_12368_48324# 0.359f
C1260 AVDD a_16040_45156# 0.356f
C1261 XA5.XA4.MN0.D a_12368_48676# 0.154f
C1262 D<2> XA6.XA3.MN0.G 0.572f
C1263 VREF XA7.XA1.XA5.MN2.D 0.341f
C1264 XA20.XA3.MN0.D XA20.XA2.MN1.D 0.617f
C1265 XA4.XA4.MN0.G XA4.XA3.MN0.G 0.554f
C1266 XA0.XA4.MN0.G XA0.XA1.XA2.MN0.D 0.206f
C1267 XA3.XA7.MN0.D a_8480_51844# 0.159f
C1268 AVDD XA8.XA4.MN0.D 2.57f
C1269 AVDD a_7328_43396# 0.361f
C1270 XA6.XA4.MN0.G a_14888_47972# 0.153f
C1271 AVDD a_5960_40932# 0.358f
C1272 AVDD a_11000_52548# 0.405f
C1273 XA3.XA3.MN0.G a_7328_45860# 0.155f
C1274 XA8.XA1.XA5.MN2.G a_18560_41636# 0.131f
C1275 AVDD XA3.XA6.MP0.G 5.93f
C1276 SARN XDAC2.X16ab.XRES1A.B 3.59f
C1277 XA0.XA1.XA5.MN2.D EN 0.162f
C1278 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES4.B 0.428f
C1279 AVDD a_12368_47268# 0.356f
C1280 SARP XA20.XA1.MN0.D 0.31f
C1281 XA0.XA7.MN0.G XA1.XA4.MN0.G 0.169f
C1282 AVDD a_12368_41636# 0.404f
C1283 SARP XDAC1.XC32a<0>.XRES1A.B 3.59f
C1284 AVDD XA0.XA11.MP0.D 0.19f
C1285 AVDD a_11000_48324# 0.359f
C1286 AVDD a_22448_42692# 0.471f
C1287 VREF XA6.XA1.XA5.MN2.D 0.341f
C1288 AVDD a_12368_54308# 0.448f
C1289 XA3.XA7.MN0.D a_7328_51844# 0.133f
C1290 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES4.B 0.428f
C1291 AVDD XA7.XA4.MN0.D 2.51f
C1292 XA6.XA1.XA5.MN2.G XA5.XA6.MP0.G 0.185f
C1293 D<2> a_16040_50788# 0.161f
C1294 AVDD a_12368_46212# 0.356f
C1295 AVDD a_5960_43396# 0.361f
C1296 XA20.XA3.MN6.D a_23600_45860# 0.154f
C1297 XB1.XA4.MN1.D a_11000_334# 0.157f
C1298 AVDD XA2.XA6.MP0.D 0.144f
C1299 CK_SAMPLE a_19928_50788# 0.164f
C1300 XA6.XA1.XA5.MN2.D a_16040_44100# 0.126f
C1301 XA20.XA2a.MN0.D XA7.XA1.XA2.MN0.D 0.227f
C1302 XA5.XA1.XA5.MN2.G D<4> 0.627f
C1303 XB1.XCAPB1.XCAPB4.A m3_7544_2420# 0.106f
C1304 AVDD a_11000_47268# 0.356f
C1305 XA7.XA6.MP0.G a_17408_50084# 0.159f
C1306 XA0.XA7.MN0.G XA0.XA4.MN0.G 0.158f
C1307 AVDD EN 40.3f
C1308 XA20.XA3a.MN0.G a_23600_46916# 0.154f
C1309 AVDD a_11000_41636# 0.404f
C1310 AVDD XA0.XA11.MN1.G 9.55f
C1311 XA1.XA10.MN0.G a_3440_52548# 0.13f
C1312 AVDD XA1.XA6.MP2.D 0.172f
C1313 XA3.XA1.XA5.MN2.D a_8480_45156# 0.153f
C1314 XA8.XA9.MN1.G XA8.XA6.MN2.D 0.126f
C1315 XDAC1.XC64b<1>.XRES2.B XDAC1.XC64b<1>.XRES16.B 0.457f
C1316 XA4.XA4.MN0.D a_11000_48676# 0.154f
C1317 AVDD a_21080_42692# 0.359f
C1318 SARP XDAC1.X16ab.XRES1A.B 3.59f
C1319 VREF XA5.XA1.XA5.MN2.D 0.341f
C1320 XA3.XA4.MN0.G XA3.XA3.MN0.G 0.639f
C1321 AVDD a_11000_54308# 0.447f
C1322 AVDD a_17408_39876# 0.438f
C1323 AVDD a_12368_51844# 0.387f
C1324 XA20.XA12.MN0.G VREF 0.188f
C1325 CK_SAMPLE a_19928_50084# 0.162f
C1326 AVDD XA6.XA4.MN0.D 2.51f
C1327 AVDD a_11000_46212# 0.356f
C1328 XA5.XA4.MN0.G a_13520_47972# 0.153f
C1329 XA20.XA3.MN6.D a_22448_45860# 0.164f
C1330 XA2.XA3.MN0.G a_5960_45860# 0.155f
C1331 XA0.XA7.MN0.G XA0.XA1.XA1.MN0.S 0.327f
C1332 CK_SAMPLE a_18560_50788# 0.157f
C1333 XDAC2.XC1.XRES8.B XDAC2.XC1.XRES2.B 0.44f
C1334 XA20.XA3a.MN0.G a_22448_46916# 0.183f
C1335 AVDD D<7> 2.23f
C1336 XA3.XA1.XA5.MN2.D a_7328_45156# 0.155f
C1337 XDAC2.XC32a<0>.XRES1A.B XDAC2.XC64a<0>.XRES1B.B 0.617f
C1338 AVDD a_12368_45156# 0.356f
C1339 XA4.XA4.MN0.D a_9848_48676# 0.158f
C1340 VREF XA4.XA1.XA5.MN2.D 0.341f
C1341 XA20.XA3.MN6.D a_22448_44804# 0.174f
C1342 AVDD a_16040_39876# 0.44f
C1343 AVDD a_11000_51844# 0.387f
C1344 DONE XA8.XA7.MN0.D 0.217f
C1345 XA2.XA7.MN0.D a_5960_51844# 0.133f
C1346 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES4.B 0.428f
C1347 CK_SAMPLE a_18560_50084# 0.167f
C1348 AVDD XA5.XA4.MN0.D 2.51f
C1349 SARN XDAC2.XC32a<0>.XRES16.B 55.3f
C1350 XA5.XA4.MN0.G a_12368_47972# 0.155f
C1351 AVDD a_2288_40932# 0.358f
C1352 AVDD a_7328_52548# 0.405f
C1353 XA2.XA3.MN0.G a_4808_45860# 0.162f
C1354 XB1.XA4.MN0.G a_9560_1038# 0.158f
C1355 AVDD XA2.XA6.MP0.G 5.93f
C1356 AVDD a_22448_44100# 0.37f
C1357 AVDD a_22448_53604# 0.37f
C1358 AVDD XA0.XA6.MP2.D 0.172f
C1359 AVDD a_7328_48324# 0.359f
C1360 AVDD a_11000_45156# 0.356f
C1361 D<3> XA5.XA3.MN0.G 0.572f
C1362 XA2.XA4.MN0.G XA2.XA3.MN0.G 0.622f
C1363 VREF XA3.XA1.XA5.MN2.D 0.341f
C1364 XA20.XA11.MN0.D DONE 0.12f
C1365 XA2.XA7.MN0.D a_4808_51844# 0.159f
C1366 AVDD XA4.XA4.MN0.D 2.51f
C1367 AVDD a_2288_43396# 0.361f
C1368 AVDD a_920_40932# 0.358f
C1369 AVDD a_5960_52548# 0.405f
C1370 XA7.XA1.XA5.MN2.G a_14888_41636# 0.128f
C1371 XA8.XA3.MN0.G a_21080_46212# 0.155f
C1372 XA0.XA11.MN1.G a_12368_2094# 0.156f
C1373 XB2.XA4.MN1.D a_12368_686# 0.161f
C1374 SARN XDAC2.X16ab.XRES16.B 55.3f
C1375 XA20.XA2a.MN0.D XA6.XA1.XA2.MN0.D 0.223f
C1376 AVDD a_7328_47268# 0.356f
C1377 XA2.XA6.MP0.G a_5960_49732# 0.101f
C1378 XDAC1.XC1.XRES8.B XDAC1.XC1.XRES2.B 0.44f
C1379 AVDD a_21080_44100# 0.359f
C1380 AVDD a_7328_41636# 0.404f
C1381 SARP XDAC1.XC32a<0>.XRES16.B 55.3f
C1382 AVDD a_21080_53604# 0.384f
C1383 AVDD a_8408_1038# 0.488f
C1384 XA2.XA1.XA5.MN2.D a_5960_45156# 0.155f
C1385 AVDD a_5960_48324# 0.359f
C1386 XA3.XA4.MN0.D a_8480_48676# 0.158f
C1387 AVDD a_17408_42692# 0.358f
C1388 VREF XA2.XA1.XA5.MN2.D 0.341f
C1389 AVDD a_7328_54308# 0.448f
C1390 AVDD XA3.XA4.MN0.D 2.65f
C1391 XDAC2.XC128a<1>.XRES8.B XDAC2.XC128a<1>.XRES2.B 0.44f
C1392 AVDD a_7328_46212# 0.356f
C1393 AVDD a_920_43396# 0.361f
C1394 XA8.XA7.MN0.G EN 0.793f
C1395 XA4.XA4.MN0.G a_11000_47972# 0.155f
C1396 XA1.XA3.MN0.G a_3440_45860# 0.162f
C1397 XA8.XA3.MN0.G a_19928_46212# 0.157f
C1398 XA0.XA11.MN1.G a_11000_2094# 0.156f
C1399 CK_SAMPLE a_14888_50788# 0.157f
C1400 AVDD XA1.XA6.MP0.D 0.144f
C1401 XA5.XA1.XA5.MN2.D a_12368_44100# 0.124f
C1402 XA4.XA1.XA5.MN2.G D<5> 0.691f
C1403 XB1.XCAPB1.XCAPB4.A m3_7544_3476# 0.106f
C1404 AVDD a_5960_47268# 0.356f
C1405 XA6.XA6.MP0.G a_16040_50084# 0.159f
C1406 AVDD a_5960_41636# 0.404f
C1407 XA0.XA10.MN0.G a_n232_52548# 0.128f
C1408 AVDD a_14960_1390# 0.434f
C1409 AVDD XA0.XA6.MP2.G 2.23f
C1410 XA2.XA1.XA5.MN2.D a_4808_45156# 0.153f
C1411 XA7.XA9.MN1.G XA7.XA6.MN2.D 0.126f
C1412 XDAC1.XC32a<0>.XRES1A.B XDAC1.XC64a<0>.XRES1B.B 0.617f
C1413 SARP a_23600_40932# 0.159f
C1414 D<3> XA3.XA3.MN0.G 0.12f
C1415 XA3.XA4.MN0.D a_7328_48676# 0.154f
C1416 AVDD a_16040_42692# 0.358f
C1417 SARP XDAC1.X16ab.XRES16.B 55.3f
C1418 XA1.XA4.MN0.G XA1.XA3.MN0.G 0.639f
C1419 VREF XA1.XA1.XA5.MN2.D 0.341f
C1420 AVDD a_5960_54308# 0.447f
C1421 AVDD a_12368_39876# 0.438f
C1422 AVDD a_7328_51844# 0.387f
C1423 XA1.XA7.MN0.D a_3440_51844# 0.159f
C1424 CK_SAMPLE a_14888_50084# 0.167f
C1425 AVDD XA2.XA4.MN0.D 2.65f
C1426 AVDD a_5960_46212# 0.356f
C1427 XA8.XA1.XA5.MN2.G EN 0.898f
C1428 XA4.XA4.MN0.G a_9848_47972# 0.153f
C1429 XA6.XA1.XA5.MN2.G a_13520_41636# 0.131f
C1430 XA1.XA3.MN0.G a_2288_45860# 0.155f
C1431 CK_SAMPLE a_13520_50788# 0.157f
C1432 AVDD XA1.XA6.MP0.G 5.92f
C1433 XDAC2.X16ab.XRES1A.B XDAC2.XC128b<2>.XRES1B.B 0.617f
C1434 XA7.XA6.MP0.G D<8> 0.132f
C1435 SARP a_23600_43396# 0.158f
C1436 AVDD a_7328_45156# 0.356f
C1437 VREF XA0.XA1.XA5.MN2.D 0.341f
C1438 XA20.XA12.MN0.G DONE 0.188f
C1439 AVDD a_11000_39876# 0.44f
C1440 AVDD a_5960_51844# 0.387f
C1441 XA1.XA7.MN0.D a_2288_51844# 0.133f
C1442 CK_SAMPLE a_13520_50084# 0.167f
C1443 AVDD XA1.XA4.MN0.D 2.65f
C1444 SARN XDAC2.XC32a<0>.XRES2.B 6.99f
C1445 D<3> a_12368_50788# 0.161f
C1446 XDAC1.XC128a<1>.XRES8.B XDAC1.XC128a<1>.XRES2.B 0.44f
C1447 AVDD XA8.XA1.XA5.MP0.D 0.143f
C1448 XA7.XA1.XA5.MN2.G EN 0.946f
C1449 AVDD a_2288_52548# 0.405f
C1450 XA7.XA3.MN0.G a_18560_46212# 0.157f
C1451 XA8.XA12.MN0.G a_19928_53604# 0.1f
C1452 AVDD XA0.XA6.MP0.D 0.144f
C1453 XA20.XA2a.MN0.D XA5.XA1.XA2.MN0.D 0.227f
C1454 XA4.XA1.XA5.MN2.D a_11000_44100# 0.126f
C1455 AVDD a_17408_44100# 0.359f
C1456 XA6.XA6.MP0.G XA2.XA3.MN0.G 0.21f
C1457 AVDD a_17408_53604# 0.383f
C1458 AVDD a_22448_51140# 0.569f
C1459 XA1.XA1.XA5.MN2.D a_3440_45156# 0.153f
C1460 XDAC2.XC64b<1>.XRES8.B XDAC2.XC64b<1>.XRES2.B 0.44f
C1461 AVDD a_2288_48324# 0.359f
C1462 AVDD a_5960_45156# 0.356f
C1463 XA2.XA4.MN0.D a_5960_48676# 0.154f
C1464 D<4> XA4.XA3.MN0.G 0.572f
C1465 XA0.XA4.MN0.G D<8> 0.622f
C1466 AVDD VREF 69.8f
C1467 XA3.XA4.MN0.G a_8480_47972# 0.153f
C1468 XA6.XA1.XA5.MN2.G EN 0.897f
C1469 AVDD a_920_52548# 0.405f
C1470 D<8> a_920_45860# 0.155f
C1471 XA7.XA3.MN0.G a_17408_46212# 0.155f
C1472 XB1.XA4.MN1.D a_11000_686# 0.161f
C1473 SARN XDAC2.X16ab.XRES2.B 6.99f
C1474 XDAC1.X16ab.XRES1A.B XDAC1.XC128b<2>.XRES1B.B 0.617f
C1475 AVDD a_2288_47268# 0.356f
C1476 AVDD a_16040_44100# 0.359f
C1477 AVDD a_2288_41636# 0.404f
C1478 SARP XDAC1.XC32a<0>.XRES2.B 6.99f
C1479 AVDD a_16040_53604# 0.383f
C1480 AVDD a_21080_51140# 0.382f
C1481 XA1.XA1.XA5.MN2.D a_2288_45156# 0.155f
C1482 AVDD a_920_48324# 0.359f
C1483 XA2.XA4.MN0.D a_4808_48676# 0.158f
C1484 D<4> XA3.XA3.MN0.G 0.225f
C1485 AVDD a_12368_42692# 0.358f
C1486 AVDD a_2288_54308# 0.448f
C1487 XA20.XA12.MN0.D XA20.XA11.MN0.D 0.178f
C1488 XA0.XA7.MN0.D a_920_51844# 0.133f
C1489 AVDD XA0.XA4.MN0.D 2.65f
C1490 XA4.XA1.XA5.MN2.G XA3.XA6.MP0.G 0.174f
C1491 XA20.XA9.MN0.D a_22448_48324# 0.139f
C1492 AVDD a_2288_46212# 0.356f
C1493 AVDD XA8.XA1.XA2.MN0.D 0.27f
C1494 XA3.XA4.MN0.G a_7328_47972# 0.155f
C1495 XA5.XA1.XA5.MN2.G EN 0.946f
C1496 D<8> a_n232_45860# 0.162f
C1497 XA7.XA12.MN0.G a_18560_53604# 0.102f
C1498 AVDD XA0.XA6.MP0.G 5.93f
C1499 CK_SAMPLE a_9848_50788# 0.157f
C1500 XA3.XA1.XA5.MN2.G D<6> 0.624f
C1501 XB2.XCAPB1.XCAPB4.A XDAC2.XC1.XRES1A.B 0.377f
C1502 XB1.XCAPB1.XCAPB4.A m3_7544_4532# 0.106f
C1503 AVDD a_920_47268# 0.356f
C1504 XA20.XA3.MN6.D XA20.XA3.MN1.D 0.159f
C1505 AVDD a_920_41636# 0.404f
C1506 XDAC1.XC64b<1>.XRES8.B XDAC1.XC64b<1>.XRES2.B 0.44f
C1507 XA8.XA4.MN0.D a_21080_49028# 0.154f
C1508 AVDD a_11000_42692# 0.358f
C1509 SARP XDAC1.X16ab.XRES2.B 6.99f
C1510 AVDD a_920_54308# 0.447f
C1511 AVDD a_7328_39876# 0.438f
C1512 AVDD a_2288_51844# 0.387f
C1513 XA8.XA7.MN0.G XA8.XA1.XA1.MP1.D 0.144f
C1514 XA20.XA3a.MN0.D EN 2.58f
C1515 XA0.XA7.MN0.D a_n232_51844# 0.159f
C1516 CK_SAMPLE a_9848_50084# 0.167f
C1517 AVDD a_920_46212# 0.356f
C1518 XA4.XA1.XA5.MN2.G EN 0.897f
C1519 AVDD XA20.XA4.MN0.D 0.456f
C1520 XA5.XA1.XA5.MN2.G a_9848_41636# 0.128f
C1521 XA6.XA3.MN0.G a_16040_46212# 0.155f
C1522 XA0.XA11.MN1.G XB2.XA4.MN1.D 0.22f
C1523 XB2.XA4.MN1.D a_12368_1038# 0.163f
C1524 XB2.XA4.MN0.G XB2.XCAPB1.XCAPB4.B 0.193f
C1525 CK_SAMPLE a_8480_50788# 0.157f
C1526 XA20.XA2a.MN0.D XA4.XA1.XA2.MN0.D 0.223f
C1527 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES8.B 0.471f
C1528 AVDD a_8408_1390# 0.435f
C1529 XA0.XA1.XA5.MN2.D a_920_45156# 0.155f
C1530 XDAC2.XC32a<0>.XRES16.B XDAC2.XC32a<0>.XRES1A.B 0.454f
C1531 AVDD a_2288_45156# 0.356f
C1532 XA1.XA4.MN0.D a_3440_48676# 0.158f
C1533 XA8.XA4.MN0.D a_19928_49028# 0.156f
C1534 AVDD a_5960_39876# 0.44f
C1535 AVDD a_920_51844# 0.387f
C1536 XA20.XA10.MN1.D XA20.XA4.MN0.D 0.11f
C1537 CK_SAMPLE a_8480_50084# 0.167f
C1538 AVDD a_22448_49732# 0.417f
C1539 SARN XDAC2.XC32a<0>.XRES8.B 27.7f
C1540 D<4> a_11000_50788# 0.161f
C1541 SARP a_23600_41636# 0.161f
C1542 D<0> XA8.XA4.MN0.G 0.239f
C1543 AVDD XA7.XA1.XA5.MP0.D 0.159f
C1544 XA2.XA4.MN0.G a_5960_47972# 0.155f
C1545 XA3.XA1.XA5.MN2.G EN 0.946f
C1546 AVDD XA8.XA10.MN0.G 0.855f
C1547 XA6.XA3.MN0.G a_14888_46212# 0.157f
C1548 XB2.XA4.MN0.G XB2.XA3.MN0.S 0.572f
C1549 AVDD a_22448_50436# 0.389f
C1550 XA3.XA1.XA5.MN2.D a_7328_44100# 0.124f
C1551 XA5.XA6.MP0.G a_12368_50084# 0.159f
C1552 XA20.XA3a.MN0.G XA20.XA3.MN6.D 1.76f
C1553 AVDD a_12368_44100# 0.359f
C1554 AVDD a_12368_53604# 0.383f
C1555 AVDD XB2.XCAPB1.XCAPB4.B 1.65f
C1556 AVDD a_17408_51140# 0.383f
C1557 XA0.XA1.XA5.MN2.D a_n232_45156# 0.153f
C1558 XA6.XA9.MN1.G XA6.XA6.MN2.D 0.126f
C1559 AVDD a_22448_48676# 0.438f
C1560 EN XA0.XA1.XA2.MN0.D 0.156f
C1561 XA8.XA7.MN0.G VREF 0.687f
C1562 AVDD a_920_45156# 0.356f
C1563 XA1.XA4.MN0.D a_2288_48676# 0.154f
C1564 D<5> XA3.XA3.MN0.G 1.2f
C1565 AVDD XA20.XA11.MP0.D 0.158f
C1566 XA20.XA12.MN0.D XA20.XA12.MN0.G 0.125f
C1567 CK_SAMPLE XA8.XA9.MN1.G 0.193f
C1568 SARN a_23600_51844# 0.156f
C1569 AVDD a_21080_49732# 0.36f
C1570 AVDD XA20.XA2a.MN0.D 9.22f
C1571 EN a_21080_42340# 0.159f
C1572 AVDD XA7.XA1.XA2.MN0.D 0.263f
C1573 XA2.XA4.MN0.G a_4808_47972# 0.153f
C1574 XA2.XA1.XA5.MN2.G EN 0.897f
C1575 XA7.XA4.MN0.G XA8.XA4.MN0.G 0.12f
C1576 AVDD XA7.XA10.MN0.G 0.853f
C1577 XA4.XA1.XA5.MN2.G a_8480_41636# 0.131f
C1578 AVDD a_21080_50436# 0.417f
C1579 SARN XDAC2.X16ab.XRES8.B 27.7f
C1580 XA20.XA2.MN1.D SARP 0.11f
C1581 AVDD a_22448_47620# 0.369f
C1582 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES8.B 0.471f
C1583 AVDD a_11000_44100# 0.359f
C1584 XA4.XA6.MP0.G XA3.XA3.MN0.G 0.271f
C1585 AVDD a_22448_41988# 0.57f
C1586 SARP XDAC1.XC32a<0>.XRES8.B 27.7f
C1587 AVDD a_11000_53604# 0.383f
C1588 AVDD XB2.XA3.MN0.S 0.183f
C1589 AVDD a_16040_51140# 0.383f
C1590 AVDD a_21080_48676# 0.356f
C1591 XA8.XA1.XA5.MN2.G VREF 0.704f
C1592 XA7.XA4.MN0.D a_18560_49028# 0.156f
C1593 AVDD a_7328_42692# 0.358f
C1594 XA8.XA7.MN0.G XA8.XA1.XA2.MN0.D 0.144f
C1595 AVDD DONE 2.49f
C1596 AVDD XA8.XA7.MN0.D 1.2f
C1597 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES8.B 0.471f
C1598 AVDD XA6.XA1.XA5.MP0.D 0.159f
C1599 XA0.XA7.MN0.G EN 0.963f
C1600 AVDD XA6.XA10.MN0.G 0.853f
C1601 XA5.XA3.MN0.G a_13520_46212# 0.157f
C1602 XA0.XA11.MN1.G XB1.XA4.MN1.D 0.216f
C1603 XB1.XA4.MN0.G XB1.XCAPB1.XCAPB4.B 0.193f
C1604 CK_SAMPLE a_4808_50788# 0.157f
C1605 XA20.XA2a.MN0.D XA3.XA1.XA2.MN0.D 0.227f
C1606 XA2.XA1.XA5.MN2.D a_5960_44100# 0.126f
C1607 XA2.XA1.XA5.MN2.G D<7> 0.691f
C1608 AVDD a_21080_47620# 0.356f
C1609 XA4.XA6.MP0.G XA2.XA3.MN0.G 0.594f
C1610 AVDD a_21080_41988# 0.386f
C1611 AVDD XB1.XCAPB1.XCAPB4.B 1.65f
C1612 XA7.XA11.MN1.G VREF 0.39f
C1613 XA7.XA1.XA5.MN2.G VREF 0.704f
C1614 XA4.XA1.XA5.MN2.G XA3.XA4.MN0.D 0.198f
C1615 XDAC1.XC32a<0>.XRES16.B XDAC1.XC32a<0>.XRES1A.B 0.454f
C1616 AVDD XA8.XA1.XA5.MN2.D 2.37f
C1617 XA7.XA4.MN0.D a_17408_49028# 0.154f
C1618 AVDD a_5960_42692# 0.358f
C1619 SARP XDAC1.X16ab.XRES8.B 27.7f
C1620 XA8.XA1.XA5.MN2.G XA8.XA1.XA2.MN0.D 0.126f
C1621 AVDD XA20.XA11.MN0.D 0.679f
C1622 AVDD a_2288_39876# 0.438f
C1623 AVDD XA7.XA7.MN0.D 1.19f
C1624 CK_SAMPLE XA7.XA9.MN1.G 0.135f
C1625 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MP1.D 0.148f
C1626 CK_SAMPLE a_4808_50084# 0.167f
C1627 AVDD a_22448_46564# 0.404f
C1628 XA1.XA4.MN0.G a_3440_47972# 0.153f
C1629 AVDD XA5.XA10.MN0.G 0.853f
C1630 XA5.XA3.MN0.G a_12368_46212# 0.155f
C1631 XA6.XA12.MN0.G a_14888_53604# 0.1f
C1632 XB1.XA4.MN1.D a_11000_1038# 0.163f
C1633 XB1.XA4.MN0.G XB1.XA3.MN0.S 0.572f
C1634 XB2.XA4.MN0.G a_14960_1742# 0.135f
C1635 CK_SAMPLE a_3440_50788# 0.157f
C1636 XB1.XCAPB1.XCAPB4.A XDAC1.XC1.XRES1A.B 0.379f
C1637 XDAC2.X16ab.XRES16.B XDAC2.X16ab.XRES1A.B 0.454f
C1638 XA0.XA6.MP0.G a_920_49732# 0.101f
C1639 XA20.XA11.MN0.D XA20.XA10.MN1.D 0.342f
C1640 AVDD XB1.XA3.MN0.S 0.183f
C1641 EN a_21080_43748# 0.166f
C1642 XA6.XA1.XA5.MN2.G VREF 0.704f
C1643 D<0> XA8.XA6.MP0.G 0.421f
C1644 AVDD XA7.XA1.XA5.MN2.D 2.36f
C1645 D<6> XA3.XA3.MN0.G 0.144f
C1646 XA0.XA4.MN0.D a_920_48676# 0.154f
C1647 AVDD a_920_39876# 0.44f
C1648 AVDD XA6.XA7.MN0.D 1.19f
C1649 AVDD a_17408_49732# 0.359f
C1650 CK_SAMPLE a_3440_50084# 0.167f
C1651 SARN XDAC2.XC32a<0>.XRES4.B 13.9f
C1652 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES8.B 0.471f
C1653 AVDD a_21080_46564# 0.356f
C1654 EN a_17408_42340# 0.159f
C1655 D<1> XA7.XA4.MN0.G 0.26f
C1656 AVDD XA6.XA1.XA2.MN0.D 0.263f
C1657 XA1.XA4.MN0.G a_2288_47972# 0.155f
C1658 AVDD XA4.XA10.MN0.G 0.853f
C1659 AVDD a_17408_50436# 0.416f
C1660 XA8.XA1.XA5.MN2.D a_21080_44452# 0.158f
C1661 XA4.XA6.MP0.G a_11000_50084# 0.159f
C1662 AVDD a_7328_44100# 0.359f
C1663 XA3.XA6.MP0.G XA3.XA3.MN0.G 3.29f
C1664 AVDD a_7328_53604# 0.383f
C1665 AVDD a_14960_1742# 0.363f
C1666 AVDD a_12368_51140# 0.383f
C1667 XA5.XA9.MN1.G XA5.XA6.MN2.D 0.126f
C1668 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES8.B 0.471f
C1669 AVDD a_17408_48676# 0.356f
C1670 XA5.XA1.XA5.MN2.G VREF 0.704f
C1671 XA3.XA1.XA5.MN2.G XA2.XA4.MN0.D 0.123f
C1672 AVDD XA6.XA1.XA5.MN2.D 2.36f
C1673 D<6> XA2.XA3.MN0.G 1.02f
C1674 XA8.XA7.MN0.G XA20.XA2a.MN0.D 0.285f
C1675 XA6.XA4.MN0.D a_16040_49028# 0.154f
C1676 XA0.XA4.MN0.D a_n232_48676# 0.158f
C1677 AVDD a_22448_54660# 0.383f
C1678 CK_SAMPLE XA6.XA9.MN1.G 0.134f
C1679 AVDD XA5.XA7.MN0.D 1.19f
C1680 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MP1.D 0.144f
C1681 AVDD a_16040_49732# 0.359f
C1682 EN a_16040_42340# 0.159f
C1683 XA5.XA4.MN0.G XA6.XA4.MN0.G 0.12f
C1684 AVDD XA3.XA10.MN0.G 0.853f
C1685 XA4.XA3.MN0.G a_11000_46212# 0.155f
C1686 XA3.XA1.XA5.MN2.G a_4808_41636# 0.128f
C1687 XA0.XA11.MN1.G a_12368_2446# 0.16f
C1688 AVDD a_16040_50436# 0.416f
C1689 SARN XDAC2.X16ab.XRES4.B 13.9f
C1690 XA20.XA2a.MN0.D XA2.XA1.XA2.MN0.D 0.223f
C1691 XA8.XA1.XA5.MN2.D a_19928_44452# 0.153f
C1692 XDAC1.X16ab.XRES16.B XDAC1.X16ab.XRES1A.B 0.454f
C1693 AVDD a_17408_47620# 0.356f
C1694 AVDD a_5960_44100# 0.359f
C1695 VREF XA20.XA3a.MN0.D 0.13f
C1696 AVDD a_17408_41988# 0.386f
C1697 SARP XDAC1.XC32a<0>.XRES4.B 13.9f
C1698 AVDD a_5960_53604# 0.383f
C1699 AVDD a_11000_51140# 0.383f
C1700 XA8.XA7.MN0.D XA8.XA7.MN0.G 0.139f
C1701 AVDD a_16040_48676# 0.356f
C1702 XA4.XA1.XA5.MN2.G VREF 0.704f
C1703 AVDD XA5.XA1.XA5.MN2.D 2.36f
C1704 XA8.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C1705 XA6.XA4.MN0.D a_14888_49028# 0.156f
C1706 AVDD a_2288_42692# 0.358f
C1707 XA8.XA1.XA5.MN2.G XA7.XA1.XA2.MN0.D 0.146f
C1708 AVDD XA20.XA12.MN0.G 1.64f
C1709 AVDD XA4.XA7.MN0.D 1.19f
C1710 D<5> a_7328_50788# 0.161f
C1711 XA2.XA1.XA5.MN2.G XA1.XA6.MP0.G 0.174f
C1712 AVDD XA5.XA1.XA5.MP0.D 0.159f
C1713 XA20.XA9.MN0.D a_23600_42692# 0.14f
C1714 XA0.XA4.MN0.G a_920_47972# 0.155f
C1715 AVDD XA2.XA10.MN0.G 0.853f
C1716 XA4.XA3.MN0.G a_9848_46212# 0.157f
C1717 XA5.XA12.MN0.G a_13520_53604# 0.102f
C1718 XA0.XA11.MN1.G a_11000_2446# 0.159f
C1719 CK_SAMPLE a_n232_50788# 0.157f
C1720 XA1.XA1.XA5.MN2.D a_2288_44100# 0.124f
C1721 XA0.XA7.MN0.G XA0.XA6.MP2.G 0.624f
C1722 AVDD a_16040_47620# 0.356f
C1723 XA8.XA7.MN0.G XA8.XA1.XA5.MN2.D 0.108f
C1724 AVDD a_16040_41988# 0.386f
C1725 XA20.XA3a.MN0.D XA8.XA1.XA2.MN0.D 0.193f
C1726 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES8.B 0.471f
C1727 XA5.XA11.MN1.G VREF 0.39f
C1728 EN a_17408_43748# 0.166f
C1729 XA3.XA1.XA5.MN2.G VREF 0.704f
C1730 XA2.XA1.XA5.MN2.G XA1.XA4.MN0.D 0.198f
C1731 AVDD XA4.XA1.XA5.MN2.D 2.36f
C1732 D<7> XA3.XA3.MN0.G 0.16f
C1733 XA7.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.51f
C1734 AVDD a_920_42692# 0.358f
C1735 SARP XDAC1.X16ab.XRES4.B 13.9f
C1736 XA7.XA1.XA5.MN2.G XA7.XA1.XA2.MN0.D 0.126f
C1737 AVDD XA20.XA12.MN0.D 1.16f
C1738 AVDD a_22448_40228# 0.47f
C1739 AVDD XA3.XA7.MN0.D 1.19f
C1740 CK_SAMPLE XA5.XA9.MN1.G 0.135f
C1741 CK_SAMPLE a_n232_50084# 0.167f
C1742 AVDD a_17408_46564# 0.356f
C1743 AVDD XA5.XA1.XA2.MN0.D 0.263f
C1744 XA0.XA4.MN0.G a_n232_47972# 0.153f
C1745 VREF XA8.XA3.MN0.G 0.603f
C1746 AVDD XA1.XA10.MN0.G 0.853f
C1747 XA2.XA1.XA5.MN2.G a_3440_41636# 0.131f
C1748 XA0.XA12.MN0.G XA0.XA11.MN1.G 0.21f
C1749 XB2.XCAPB1.XCAPB4.A XB2.XCAPB1.XCAPB4.B 0.376p
C1750 XA7.XA1.XA5.MN2.D a_18560_44452# 0.153f
C1751 EN a_21080_43044# 0.14f
C1752 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES4.B 0.428f
C1753 XA2.XA6.MP0.G XA3.XA3.MN0.G 3.56f
C1754 XA20.XA12.MN0.G XA8.XA12.MN0.G 0.124f
C1755 XA20.XA12.MN0.D XA20.XA10.MN1.D 0.125f
C1756 XA7.XA7.MN0.D XA8.XA1.XA5.MN2.G 0.14f
C1757 EN a_16040_43748# 0.166f
C1758 XA2.XA1.XA5.MN2.G VREF 0.704f
C1759 AVDD XA3.XA1.XA5.MN2.D 2.36f
C1760 D<7> XA2.XA3.MN0.G 0.112f
C1761 XA6.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C1762 XA5.XA4.MN0.D a_13520_49028# 0.156f
C1763 AVDD a_21080_40228# 0.469f
C1764 AVDD XA2.XA7.MN0.D 1.19f
C1765 AVDD a_12368_49732# 0.359f
C1766 SARN XDAC2.XC32a<0>.XRES1B.B 3.59f
C1767 AVDD a_16040_46564# 0.356f
C1768 EN a_12368_42340# 0.159f
C1769 D<2> XA6.XA4.MN0.G 0.26f
C1770 AVDD XA4.XA1.XA5.MP0.D 0.159f
C1771 XA20.XA3.MN0.D XA20.XA2a.MN0.D 0.218f
C1772 VREF XA7.XA3.MN0.G 0.608f
C1773 AVDD XA0.XA10.MN0.G 0.853f
C1774 XA3.XA3.MN0.G a_8480_46212# 0.157f
C1775 AVDD a_12368_50436# 0.416f
C1776 XA20.XA2a.MN0.D XA1.XA1.XA2.MN0.D 0.227f
C1777 XA0.XA1.XA5.MN2.D a_920_44100# 0.126f
C1778 XA7.XA1.XA5.MN2.D a_17408_44452# 0.158f
C1779 AVDD a_2288_44100# 0.359f
C1780 XA2.XA6.MP0.G XA2.XA3.MN0.G 3.15f
C1781 XA8.XA1.XA5.MN2.G XA7.XA1.XA5.MN2.D 0.108f
C1782 AVDD a_2288_53604# 0.383f
C1783 AVDD a_7328_51140# 0.383f
C1784 D<8> EN 0.298f
C1785 AVDD a_12368_48676# 0.356f
C1786 XA0.XA7.MN0.G VREF 0.704f
C1787 XDAC2.XC32a<0>.XRES2.B XDAC2.XC32a<0>.XRES16.B 0.457f
C1788 AVDD XA2.XA1.XA5.MN2.D 2.36f
C1789 D<7> XA1.XA3.MN0.G 1.21f
C1790 XA5.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.51f
C1791 XA5.XA4.MN0.D a_12368_49028# 0.154f
C1792 AVDD a_22448_55012# 0.467f
C1793 AVDD XA1.XA7.MN0.D 1.19f
C1794 CK_SAMPLE XA4.XA9.MN1.G 0.134f
C1795 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MP1.D 0.148f
C1796 AVDD a_11000_49732# 0.359f
C1797 D<2> D<1> 6.86f
C1798 XB2.XCAPB1.XCAPB4.B m3_26048_132# 0.17f
C1799 EN a_11000_42340# 0.159f
C1800 XA3.XA4.MN0.D XA3.XA3.MN0.G 0.158f
C1801 XA3.XA4.MN0.G XA4.XA4.MN0.G 0.12f
C1802 VREF XA6.XA3.MN0.G 0.608f
C1803 XA3.XA3.MN0.G a_7328_46212# 0.155f
C1804 XB1.XA4.MN0.G a_8408_1742# 0.135f
C1805 AVDD a_11000_50436# 0.416f
C1806 SARN XDAC2.X16ab.XRES1B.B 3.59f
C1807 AVDD a_12368_47620# 0.356f
C1808 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES4.B 0.428f
C1809 AVDD a_920_44100# 0.359f
C1810 AVDD a_12368_41988# 0.386f
C1811 SARP XDAC1.XC32a<0>.XRES1B.B 3.59f
C1812 XA20.XA3a.MN0.D XA20.XA2a.MN0.D 3.6f
C1813 AVDD a_920_53604# 0.383f
C1814 AVDD a_8408_1742# 0.363f
C1815 AVDD a_5960_51140# 0.383f
C1816 XA0.XA11.MN1.G SARN 0.393f
C1817 XA20.XA3a.MN0.D XA7.XA1.XA2.MN0.D 0.199f
C1818 XA6.XA7.MN0.D XA7.XA1.XA5.MN2.G 0.14f
C1819 AVDD a_11000_48676# 0.356f
C1820 XA0.XA7.MN0.G XA0.XA4.MN0.D 0.123f
C1821 D<1> XA7.XA6.MP0.G 3.47f
C1822 AVDD XA1.XA1.XA5.MN2.D 2.36f
C1823 XA0.XA6.MP2.G XA3.XA3.MN0.G 0.347f
C1824 XA4.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C1825 XA7.XA1.XA5.MN2.G XA6.XA1.XA2.MN0.D 0.144f
C1826 AVDD XA0.XA7.MN0.D 1.19f
C1827 D<6> a_5960_50788# 0.161f
C1828 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES4.B 0.428f
C1829 XA0.XA11.MN1.G SARP 0.523f
C1830 AVDD XA4.XA1.XA2.MN0.D 0.263f
C1831 XA2.XA4.MN0.D XA3.XA3.MN0.G 0.11f
C1832 XA20.XA3.MN6.D a_23600_46212# 0.154f
C1833 VREF XA5.XA3.MN0.G 0.608f
C1834 AVDD a_22448_52900# 0.486f
C1835 XA0.XA11.MN1.G SAR_IN 0.377f
C1836 XA6.XA1.XA5.MN2.D a_16040_44452# 0.158f
C1837 AVDD a_11000_47620# 0.356f
C1838 EN a_17408_43044# 0.141f
C1839 XA3.XA6.MP0.G a_7328_50084# 0.159f
C1840 XA20.XA3a.MN0.G a_23600_47268# 0.154f
C1841 XA1.XA6.MP0.G XA3.XA3.MN0.G 0.214f
C1842 XA7.XA1.XA5.MN2.G XA6.XA1.XA5.MN2.D 0.108f
C1843 AVDD a_11000_41988# 0.386f
C1844 AVDD XB2.XA4.MN0.G 2.28f
C1845 XA4.XA9.MN1.G XA4.XA6.MN2.D 0.126f
C1846 XA3.XA11.MN1.G VREF 0.39f
C1847 SARN XDAC2.XC1.XRES1A.B 3.59f
C1848 EN a_12368_43748# 0.166f
C1849 XDAC1.XC32a<0>.XRES2.B XDAC1.XC32a<0>.XRES16.B 0.457f
C1850 AVDD XA0.XA1.XA5.MN2.D 2.36f
C1851 XA0.XA6.MP2.G XA2.XA3.MN0.G 0.675f
C1852 XA3.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.51f
C1853 XA4.XA4.MN0.D a_11000_49028# 0.154f
C1854 SARP XDAC1.X16ab.XRES1B.B 3.59f
C1855 XA6.XA1.XA5.MN2.G XA6.XA1.XA2.MN0.D 0.126f
C1856 AVDD a_22448_55364# 0.448f
C1857 AVDD a_17408_40228# 0.464f
C1858 CK_SAMPLE XA3.XA9.MN1.G 0.135f
C1859 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MP1.D 0.144f
C1860 SARP a_23600_44100# 0.154f
C1861 AVDD a_12368_46564# 0.356f
C1862 XA1.XA4.MN0.D XA3.XA3.MN0.G 0.113f
C1863 D<7> SARP 0.137f
C1864 XA20.XA3.MN6.D a_22448_46212# 0.164f
C1865 VREF XA4.XA3.MN0.G 0.608f
C1866 AVDD a_21080_52900# 0.387f
C1867 XA2.XA3.MN0.G a_5960_46212# 0.155f
C1868 XA0.XA7.MN0.G a_n232_41636# 0.128f
C1869 XA4.XA12.MN0.G a_9848_53604# 0.1f
C1870 XA20.XA2a.MN0.D XA0.XA1.XA2.MN0.D 0.223f
C1871 XA6.XA1.XA5.MN2.D a_14888_44452# 0.153f
C1872 XDAC2.X16ab.XRES2.B XDAC2.X16ab.XRES16.B 0.457f
C1873 EN a_16040_43044# 0.141f
C1874 XA20.XA3a.MN0.G a_22448_47268# 0.182f
C1875 XA1.XA6.MP0.G XA2.XA3.MN0.G 5.91f
C1876 AVDD XB1.XA4.MN0.G 2.28f
C1877 XA5.XA7.MN0.D XA6.XA1.XA5.MN2.G 0.14f
C1878 EN a_11000_43748# 0.166f
C1879 XA0.XA6.MP2.G XA1.XA3.MN0.G 0.194f
C1880 XA2.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C1881 XA4.XA4.MN0.D a_9848_49028# 0.156f
C1882 XA8.XA4.MN0.G a_21080_47268# 0.155f
C1883 XA20.XA3a.MN0.G XA20.XA2.MN1.D 0.126f
C1884 XA20.XA3.MN6.D a_23600_45156# 0.134f
C1885 AVDD a_16040_40228# 0.467f
C1886 AVDD a_22448_52196# 0.569f
C1887 AVDD a_7328_49732# 0.359f
C1888 SARN XDAC2.XC128a<1>.XRES1A.B 3.59f
C1889 D<3> D<1> 0.356f
C1890 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES4.B 0.428f
C1891 AVDD a_11000_46564# 0.356f
C1892 EN a_7328_42340# 0.159f
C1893 D<3> XA5.XA4.MN0.G 0.26f
C1894 AVDD XA3.XA1.XA5.MP0.D 0.159f
C1895 XA1.XA4.MN0.D XA2.XA3.MN0.G 0.109f
C1896 VREF XA3.XA3.MN0.G 0.608f
C1897 SARP XDAC1.XC1.XRES1A.B 3.59f
C1898 XA2.XA3.MN0.G a_4808_46212# 0.157f
C1899 XA20.XA10.MN1.D XA20.XA10.MN0.D 0.142f
C1900 XA0.XA11.MN1.G SAR_IP 0.374f
C1901 AVDD a_7328_50436# 0.416f
C1902 AVDD a_22448_44452# 0.416f
C1903 XA6.XA1.XA5.MN2.G XA5.XA1.XA5.MN2.D 0.108f
C1904 XA1.XA6.MP0.G XA1.XA3.MN0.G 2.44f
C1905 AVDD XA20.XA10.MN1.D 2.12f
C1906 AVDD a_14960_2094# 0.362f
C1907 AVDD a_2288_51140# 0.383f
C1908 XA20.XA3a.MN0.D XA6.XA1.XA2.MN0.D 0.195f
C1909 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES4.B 0.428f
C1910 AVDD a_7328_48676# 0.356f
C1911 D<2> XA7.XA6.MP0.G 0.112f
C1912 AVDD a_22448_45508# 0.368f
C1913 EN XA8.XA1.XA1.MN0.S 0.139f
C1914 XA0.XA6.MP2.G D<8> 1.31f
C1915 XA0.XA7.MN0.G XA20.XA2a.MN0.D 0.51f
C1916 XA8.XA4.MN0.G a_19928_47268# 0.157f
C1917 XA20.XA3.MN6.D a_22448_45156# 0.15f
C1918 AVDD a_21080_52196# 0.37f
C1919 CK_SAMPLE XA2.XA9.MN1.G 0.134f
C1920 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D 0.702f
C1921 AVDD a_5960_49732# 0.359f
C1922 XB2.XCAPB1.XCAPB4.B m3_26048_1188# 0.17f
C1923 EN a_5960_42340# 0.159f
C1924 AVDD XA3.XA1.XA2.MN0.D 0.263f
C1925 XA1.XA4.MN0.G XA2.XA4.MN0.G 0.12f
C1926 VREF XA2.XA3.MN0.G 0.608f
C1927 XA0.XA4.MN0.D XA3.XA3.MN0.G 0.123f
C1928 XA1.XA4.MN0.D XA1.XA3.MN0.G 0.157f
C1929 XB1.XCAPB1.XCAPB4.A XB1.XCAPB1.XCAPB4.B 0.376p
C1930 AVDD a_5960_50436# 0.416f
C1931 XA5.XA1.XA5.MN2.D a_13520_44452# 0.153f
C1932 SARN XDAC2.XC64b<1>.XRES1A.B 3.59f
C1933 XDAC1.X16ab.XRES2.B XDAC1.X16ab.XRES16.B 0.457f
C1934 AVDD a_7328_47620# 0.356f
C1935 AVDD a_21080_44452# 0.357f
C1936 XA0.XA6.MP0.G XA3.XA3.MN0.G 0.326f
C1937 AVDD a_7328_41988# 0.386f
C1938 SARP XDAC1.XC128a<1>.XRES1A.B 3.59f
C1939 AVDD XA8.XA12.MN0.G 0.71f
C1940 AVDD a_920_51140# 0.383f
C1941 XA4.XA7.MN0.D XA5.XA1.XA5.MN2.G 0.14f
C1942 AVDD a_5960_48676# 0.356f
C1943 AVDD a_21080_45508# 0.359f
C1944 XA3.XA4.MN0.D a_8480_49028# 0.156f
C1945 XA6.XA1.XA5.MN2.G XA5.XA1.XA2.MN0.D 0.146f
C1946 AVDD XA2.XA1.XA5.MP0.D 0.159f
C1947 VREF XA1.XA3.MN0.G 0.608f
C1948 XA0.XA4.MN0.D XA2.XA3.MN0.G 0.11f
C1949 XA0.XA6.MP2.G SARP 0.312f
C1950 AVDD a_22448_41284# 0.569f
C1951 AVDD a_17408_52900# 0.387f
C1952 XA1.XA3.MN0.G a_3440_46212# 0.157f
C1953 XA8.XA3.MN0.G a_21080_46564# 0.155f
C1954 XA3.XA12.MN0.G a_8480_53604# 0.102f
C1955 XA5.XA1.XA5.MN2.D a_12368_44452# 0.158f
C1956 SARN XA1.XA6.MP0.G 0.171f
C1957 AVDD a_5960_47620# 0.356f
C1958 EN a_12368_43044# 0.141f
C1959 XA2.XA6.MP0.G a_5960_50084# 0.159f
C1960 XA5.XA1.XA5.MN2.G XA4.XA1.XA5.MN2.D 0.108f
C1961 XA0.XA6.MP0.G XA2.XA3.MN0.G 0.133f
C1962 AVDD a_5960_41988# 0.386f
C1963 AVDD XA7.XA12.MN0.G 0.706f
C1964 XDAC2.XC1.XRES1A.B AVSS 8.27f
C1965 XDAC1.XC1.XRES1A.B AVSS 8.27f
C1966 XDAC2.XC1.XRES16.B AVSS 22.8f
C1967 XDAC1.XC1.XRES16.B AVSS 22.8f
C1968 XDAC2.XC1.XRES2.B AVSS 9.09f
C1969 XDAC1.XC1.XRES2.B AVSS 9.09f
C1970 XDAC2.XC1.XRES8.B AVSS 15f
C1971 XDAC1.XC1.XRES8.B AVSS 15f
C1972 XDAC2.XC1.XRES4.B AVSS 11.1f
C1973 XDAC1.XC1.XRES4.B AVSS 11.1f
C1974 XDAC2.XC1.XRES1B.B AVSS 8.07f
C1975 XDAC1.XC1.XRES1B.B AVSS 8.07f
C1976 XDAC2.XC64a<0>.XRES1A.B AVSS 8.06f
C1977 XDAC1.XC64a<0>.XRES1A.B AVSS 8.06f
C1978 XDAC2.XC64a<0>.XRES16.B AVSS 22.8f
C1979 XDAC1.XC64a<0>.XRES16.B AVSS 22.8f
C1980 XDAC2.XC64a<0>.XRES2.B AVSS 9.09f
C1981 XDAC1.XC64a<0>.XRES2.B AVSS 9.09f
C1982 XDAC2.XC64a<0>.XRES8.B AVSS 15f
C1983 XDAC1.XC64a<0>.XRES8.B AVSS 15f
C1984 XDAC2.XC64a<0>.XRES4.B AVSS 11.1f
C1985 XDAC1.XC64a<0>.XRES4.B AVSS 11.1f
C1986 XDAC2.XC64a<0>.XRES1B.B AVSS 8.07f
C1987 XDAC1.XC64a<0>.XRES1B.B AVSS 8.07f
C1988 XDAC2.XC32a<0>.XRES1A.B AVSS 8.06f
C1989 XDAC1.XC32a<0>.XRES1A.B AVSS 8.06f
C1990 XDAC2.XC32a<0>.XRES16.B AVSS 22.8f
C1991 XDAC1.XC32a<0>.XRES16.B AVSS 22.8f
C1992 XDAC2.XC32a<0>.XRES2.B AVSS 9.09f
C1993 XDAC1.XC32a<0>.XRES2.B AVSS 9.09f
C1994 XDAC2.XC32a<0>.XRES8.B AVSS 15f
C1995 XDAC1.XC32a<0>.XRES8.B AVSS 15f
C1996 XDAC2.XC32a<0>.XRES4.B AVSS 11.1f
C1997 XDAC1.XC32a<0>.XRES4.B AVSS 11.1f
C1998 XDAC2.XC32a<0>.XRES1B.B AVSS 8.07f
C1999 XDAC1.XC32a<0>.XRES1B.B AVSS 8.07f
C2000 XDAC2.XC128a<1>.XRES1A.B AVSS 8.06f
C2001 XDAC1.XC128a<1>.XRES1A.B AVSS 8.06f
C2002 XDAC2.XC128a<1>.XRES16.B AVSS 22.8f
C2003 XDAC1.XC128a<1>.XRES16.B AVSS 22.8f
C2004 XDAC2.XC128a<1>.XRES2.B AVSS 9.09f
C2005 XDAC1.XC128a<1>.XRES2.B AVSS 9.09f
C2006 XDAC2.XC128a<1>.XRES8.B AVSS 15f
C2007 XDAC1.XC128a<1>.XRES8.B AVSS 15f
C2008 XDAC2.XC128a<1>.XRES4.B AVSS 11.1f
C2009 XDAC1.XC128a<1>.XRES4.B AVSS 11.1f
C2010 XDAC2.XC128a<1>.XRES1B.B AVSS 8.07f
C2011 XDAC1.XC128a<1>.XRES1B.B AVSS 8.07f
C2012 XDAC2.XC128b<2>.XRES1A.B AVSS 8.06f
C2013 XDAC1.XC128b<2>.XRES1A.B AVSS 8.06f
C2014 XDAC2.XC128b<2>.XRES16.B AVSS 22.8f
C2015 XDAC1.XC128b<2>.XRES16.B AVSS 22.8f
C2016 XDAC2.XC128b<2>.XRES2.B AVSS 9.09f
C2017 XDAC1.XC128b<2>.XRES2.B AVSS 9.09f
C2018 XDAC2.XC128b<2>.XRES8.B AVSS 15f
C2019 XDAC1.XC128b<2>.XRES8.B AVSS 15f
C2020 XDAC2.XC128b<2>.XRES4.B AVSS 11.1f
C2021 XDAC1.XC128b<2>.XRES4.B AVSS 11.1f
C2022 XDAC2.XC128b<2>.XRES1B.B AVSS 8.07f
C2023 XDAC1.XC128b<2>.XRES1B.B AVSS 8.07f
C2024 XDAC2.X16ab.XRES1A.B AVSS 8.06f
C2025 XDAC1.X16ab.XRES1A.B AVSS 8.06f
C2026 XDAC2.X16ab.XRES16.B AVSS 22.8f
C2027 XDAC1.X16ab.XRES16.B AVSS 22.8f
C2028 XDAC2.X16ab.XRES2.B AVSS 9.09f
C2029 XDAC1.X16ab.XRES2.B AVSS 9.09f
C2030 XDAC2.X16ab.XRES8.B AVSS 15f
C2031 XDAC1.X16ab.XRES8.B AVSS 15f
C2032 XDAC2.X16ab.XRES4.B AVSS 11.1f
C2033 XDAC1.X16ab.XRES4.B AVSS 11.1f
C2034 XDAC2.X16ab.XRES1B.B AVSS 8.07f
C2035 XDAC1.X16ab.XRES1B.B AVSS 8.07f
C2036 XDAC2.XC64b<1>.XRES1A.B AVSS 8.06f
C2037 XDAC1.XC64b<1>.XRES1A.B AVSS 8.06f
C2038 XDAC2.XC64b<1>.XRES16.B AVSS 22.8f
C2039 XDAC1.XC64b<1>.XRES16.B AVSS 22.8f
C2040 XDAC2.XC64b<1>.XRES2.B AVSS 9.09f
C2041 XDAC1.XC64b<1>.XRES2.B AVSS 9.09f
C2042 XDAC2.XC64b<1>.XRES8.B AVSS 15f
C2043 XDAC1.XC64b<1>.XRES8.B AVSS 15f
C2044 XDAC2.XC64b<1>.XRES4.B AVSS 11.1f
C2045 XDAC1.XC64b<1>.XRES4.B AVSS 11.1f
C2046 XDAC2.XC64b<1>.XRES1B.B AVSS 8.07f
C2047 XDAC1.XC64b<1>.XRES1B.B AVSS 8.07f
C2048 XDAC2.XC0.XRES1A.B AVSS 8.06f
C2049 XDAC1.XC0.XRES1A.B AVSS 8.06f
C2050 XDAC2.XC0.XRES16.B AVSS 22.8f
C2051 XDAC1.XC0.XRES16.B AVSS 22.8f
C2052 XDAC2.XC0.XRES2.B AVSS 9.09f
C2053 XDAC1.XC0.XRES2.B AVSS 9.09f
C2054 XDAC2.XC0.XRES8.B AVSS 15f
C2055 XDAC1.XC0.XRES8.B AVSS 15f
C2056 XDAC2.XC0.XRES4.B AVSS 11.1f
C2057 XDAC1.XC0.XRES4.B AVSS 11.1f
C2058 XDAC2.XC0.XRES1B.B AVSS 8.75f
C2059 XDAC1.XC0.XRES1B.B AVSS 8.75f
C2060 a_13808_n18# AVSS 0.539f $ **FLOATING
C2061 a_12368_n18# AVSS 0.428f $ **FLOATING
C2062 a_11000_n18# AVSS 0.427f $ **FLOATING
C2063 a_9560_n18# AVSS 0.54f $ **FLOATING
C2064 a_13808_334# AVSS 0.488f $ **FLOATING
C2065 a_12368_334# AVSS 0.353f $ **FLOATING
C2066 a_11000_334# AVSS 0.353f $ **FLOATING
C2067 a_9560_334# AVSS 0.487f $ **FLOATING
C2068 CK_SAMPLE_BSSW AVSS 28.3f
C2069 a_13808_686# AVSS 0.365f $ **FLOATING
C2070 a_12368_686# AVSS 0.352f $ **FLOATING
C2071 a_11000_686# AVSS 0.352f $ **FLOATING
C2072 a_9560_686# AVSS 0.365f $ **FLOATING
C2073 a_13808_1038# AVSS 0.414f $ **FLOATING
C2074 a_12368_1038# AVSS 0.352f $ **FLOATING
C2075 a_11000_1038# AVSS 0.352f $ **FLOATING
C2076 a_9560_1038# AVSS 0.414f $ **FLOATING
C2077 a_13808_1390# AVSS 0.363f $ **FLOATING
C2078 a_12368_1390# AVSS 0.354f $ **FLOATING
C2079 a_11000_1390# AVSS 0.354f $ **FLOATING
C2080 a_9560_1390# AVSS 0.363f $ **FLOATING
C2081 XB2.XCAPB1.XCAPB4.B AVSS 52.2f
C2082 XB2.XA3.MN0.S AVSS 0.813f
C2083 XB1.XCAPB1.XCAPB4.B AVSS 52.2f
C2084 XB1.XA3.MN0.S AVSS 0.813f
C2085 a_13808_1742# AVSS 0.382f $ **FLOATING
C2086 a_12368_1742# AVSS 0.352f $ **FLOATING
C2087 a_11000_1742# AVSS 0.352f $ **FLOATING
C2088 a_9560_1742# AVSS 0.382f $ **FLOATING
C2089 XB2.XA4.MN0.G AVSS 2.63f
C2090 XB1.XA4.MN0.G AVSS 2.63f
C2091 a_13808_2094# AVSS 0.363f $ **FLOATING
C2092 a_12368_2094# AVSS 0.352f $ **FLOATING
C2093 a_11000_2094# AVSS 0.352f $ **FLOATING
C2094 a_9560_2094# AVSS 0.363f $ **FLOATING
C2095 XB2.XCAPB1.XCAPB4.A AVSS 49f
C2096 XB2.XA4.MN0.D AVSS 0.162f
C2097 XB2.XA4.MN1.D AVSS 3.18f
C2098 XB1.XA4.MN0.D AVSS 0.162f
C2099 XB1.XCAPB1.XCAPB4.A AVSS 49f
C2100 XB1.XA4.MN1.D AVSS 3.12f
C2101 a_13808_2446# AVSS 0.382f $ **FLOATING
C2102 a_12368_2446# AVSS 0.352f $ **FLOATING
C2103 a_11000_2446# AVSS 0.352f $ **FLOATING
C2104 a_9560_2446# AVSS 0.382f $ **FLOATING
C2105 XB2.XA4.MN1.G AVSS 0.941f
C2106 SAR_IN AVSS 1.81f
C2107 XB2.XA1.MN0.D AVSS 0.786f
C2108 SAR_IP AVSS 1.81f
C2109 XB1.XA1.MN0.D AVSS 0.786f
C2110 XB1.XA4.MN1.G AVSS 0.941f
C2111 a_13808_2798# AVSS 0.467f $ **FLOATING
C2112 a_12368_2798# AVSS 0.422f $ **FLOATING
C2113 a_11000_2798# AVSS 0.423f $ **FLOATING
C2114 a_9560_2798# AVSS 0.468f $ **FLOATING
C2115 a_13808_3150# AVSS 0.49f $ **FLOATING
C2116 XB2.XA2.MN0.G AVSS 0.591f
C2117 a_13808_3502# AVSS 0.468f $ **FLOATING
C2118 a_13808_3854# AVSS 0.538f $ **FLOATING
C2119 a_9560_3150# AVSS 0.489f $ **FLOATING
C2120 XB1.XA2.MN0.G AVSS 0.591f
C2121 a_9560_3502# AVSS 0.47f $ **FLOATING
C2122 a_9560_3854# AVSS 0.537f $ **FLOATING
C2123 a_23600_39876# AVSS 0.529f $ **FLOATING
C2124 a_19928_39876# AVSS 0.528f $ **FLOATING
C2125 a_18560_39876# AVSS 0.529f $ **FLOATING
C2126 a_14888_39876# AVSS 0.528f $ **FLOATING
C2127 a_13520_39876# AVSS 0.529f $ **FLOATING
C2128 a_9848_39876# AVSS 0.527f $ **FLOATING
C2129 a_8480_39876# AVSS 0.528f $ **FLOATING
C2130 a_4808_39876# AVSS 0.527f $ **FLOATING
C2131 a_3440_39876# AVSS 0.528f $ **FLOATING
C2132 a_n232_39876# AVSS 0.528f $ **FLOATING
C2133 a_23600_40228# AVSS 0.487f $ **FLOATING
C2134 a_19928_40228# AVSS 0.469f $ **FLOATING
C2135 a_18560_40228# AVSS 0.463f $ **FLOATING
C2136 a_14888_40228# AVSS 0.469f $ **FLOATING
C2137 a_13520_40228# AVSS 0.463f $ **FLOATING
C2138 a_9848_40228# AVSS 0.468f $ **FLOATING
C2139 a_8480_40228# AVSS 0.461f $ **FLOATING
C2140 a_4808_40228# AVSS 0.468f $ **FLOATING
C2141 a_3440_40228# AVSS 0.461f $ **FLOATING
C2142 a_n232_40228# AVSS 0.469f $ **FLOATING
C2143 a_23600_40580# AVSS 0.363f $ **FLOATING
C2144 a_19928_40580# AVSS 0.385f $ **FLOATING
C2145 a_18560_40580# AVSS 0.384f $ **FLOATING
C2146 a_14888_40580# AVSS 0.385f $ **FLOATING
C2147 a_13520_40580# AVSS 0.384f $ **FLOATING
C2148 a_9848_40580# AVSS 0.385f $ **FLOATING
C2149 a_8480_40580# AVSS 0.382f $ **FLOATING
C2150 a_4808_40580# AVSS 0.384f $ **FLOATING
C2151 a_3440_40580# AVSS 0.382f $ **FLOATING
C2152 a_n232_40580# AVSS 0.385f $ **FLOATING
C2153 a_23600_40932# AVSS 0.358f $ **FLOATING
C2154 a_19928_40932# AVSS 0.369f $ **FLOATING
C2155 a_18560_40932# AVSS 0.367f $ **FLOATING
C2156 a_14888_40932# AVSS 0.369f $ **FLOATING
C2157 a_13520_40932# AVSS 0.367f $ **FLOATING
C2158 a_9848_40932# AVSS 0.368f $ **FLOATING
C2159 a_8480_40932# AVSS 0.366f $ **FLOATING
C2160 a_4808_40932# AVSS 0.368f $ **FLOATING
C2161 a_3440_40932# AVSS 0.366f $ **FLOATING
C2162 a_n232_40932# AVSS 0.369f $ **FLOATING
C2163 XA8.XA1.XA1.MN0.D AVSS 0.478f
C2164 XA7.XA1.XA1.MN0.D AVSS 0.451f
C2165 XA6.XA1.XA1.MN0.D AVSS 0.474f
C2166 XA5.XA1.XA1.MN0.D AVSS 0.451f
C2167 XA4.XA1.XA1.MN0.D AVSS 0.474f
C2168 XA3.XA1.XA1.MN0.D AVSS 0.451f
C2169 XA2.XA1.XA1.MN0.D AVSS 0.474f
C2170 XA1.XA1.XA1.MN0.D AVSS 0.451f
C2171 XA0.XA1.XA1.MN0.D AVSS 0.474f
C2172 a_23600_41284# AVSS 0.357f $ **FLOATING
C2173 a_19928_41284# AVSS 0.404f $ **FLOATING
C2174 a_18560_41284# AVSS 0.404f $ **FLOATING
C2175 a_14888_41284# AVSS 0.404f $ **FLOATING
C2176 a_13520_41284# AVSS 0.404f $ **FLOATING
C2177 a_9848_41284# AVSS 0.403f $ **FLOATING
C2178 a_8480_41284# AVSS 0.402f $ **FLOATING
C2179 a_4808_41284# AVSS 0.403f $ **FLOATING
C2180 a_3440_41284# AVSS 0.402f $ **FLOATING
C2181 a_n232_41284# AVSS 0.404f $ **FLOATING
C2182 XA8.XA1.XA1.MN0.S AVSS 0.745f
C2183 XA7.XA1.XA1.MN0.S AVSS 0.728f
C2184 XA6.XA1.XA1.MN0.S AVSS 0.738f
C2185 XA5.XA1.XA1.MN0.S AVSS 0.728f
C2186 XA4.XA1.XA1.MN0.S AVSS 0.737f
C2187 XA3.XA1.XA1.MN0.S AVSS 0.725f
C2188 XA2.XA1.XA1.MN0.S AVSS 0.736f
C2189 XA1.XA1.XA1.MN0.S AVSS 0.724f
C2190 XA0.XA1.XA1.MN0.S AVSS 0.738f
C2191 a_23600_41636# AVSS 0.357f $ **FLOATING
C2192 a_19928_41636# AVSS 0.386f $ **FLOATING
C2193 a_18560_41636# AVSS 0.386f $ **FLOATING
C2194 a_14888_41636# AVSS 0.386f $ **FLOATING
C2195 a_13520_41636# AVSS 0.386f $ **FLOATING
C2196 a_9848_41636# AVSS 0.385f $ **FLOATING
C2197 a_8480_41636# AVSS 0.384f $ **FLOATING
C2198 a_4808_41636# AVSS 0.385f $ **FLOATING
C2199 a_3440_41636# AVSS 0.384f $ **FLOATING
C2200 a_n232_41636# AVSS 0.386f $ **FLOATING
C2201 a_23600_41988# AVSS 0.357f $ **FLOATING
C2202 a_19928_41988# AVSS 0.385f $ **FLOATING
C2203 a_18560_41988# AVSS 0.386f $ **FLOATING
C2204 a_14888_41988# AVSS 0.386f $ **FLOATING
C2205 a_13520_41988# AVSS 0.386f $ **FLOATING
C2206 a_9848_41988# AVSS 0.385f $ **FLOATING
C2207 a_8480_41988# AVSS 0.384f $ **FLOATING
C2208 a_4808_41988# AVSS 0.385f $ **FLOATING
C2209 a_3440_41988# AVSS 0.384f $ **FLOATING
C2210 a_n232_41988# AVSS 0.386f $ **FLOATING
C2211 a_23600_42340# AVSS 0.36f $ **FLOATING
C2212 a_19928_42340# AVSS 0.36f $ **FLOATING
C2213 a_18560_42340# AVSS 0.36f $ **FLOATING
C2214 a_14888_42340# AVSS 0.361f $ **FLOATING
C2215 a_13520_42340# AVSS 0.36f $ **FLOATING
C2216 a_9848_42340# AVSS 0.36f $ **FLOATING
C2217 a_8480_42340# AVSS 0.359f $ **FLOATING
C2218 a_4808_42340# AVSS 0.36f $ **FLOATING
C2219 a_3440_42340# AVSS 0.359f $ **FLOATING
C2220 a_n232_42340# AVSS 0.361f $ **FLOATING
C2221 XA20.XA1.MN0.D AVSS 0.946f
C2222 XA8.XA1.XA4.MN0.D AVSS 0.134f
C2223 XA7.XA1.XA4.MN0.D AVSS 0.139f
C2224 XA6.XA1.XA4.MN0.D AVSS 0.139f
C2225 XA5.XA1.XA4.MN0.D AVSS 0.139f
C2226 XA4.XA1.XA4.MN0.D AVSS 0.139f
C2227 XA3.XA1.XA4.MN0.D AVSS 0.139f
C2228 XA2.XA1.XA4.MN0.D AVSS 0.139f
C2229 XA1.XA1.XA4.MN0.D AVSS 0.139f
C2230 XA0.XA1.XA4.MN0.D AVSS 0.139f
C2231 a_23600_42692# AVSS 0.381f $ **FLOATING
C2232 a_19928_42692# AVSS 0.358f $ **FLOATING
C2233 a_18560_42692# AVSS 0.357f $ **FLOATING
C2234 a_14888_42692# AVSS 0.357f $ **FLOATING
C2235 a_13520_42692# AVSS 0.357f $ **FLOATING
C2236 a_9848_42692# AVSS 0.356f $ **FLOATING
C2237 a_8480_42692# AVSS 0.355f $ **FLOATING
C2238 a_4808_42692# AVSS 0.356f $ **FLOATING
C2239 a_3440_42692# AVSS 0.355f $ **FLOATING
C2240 a_n232_42692# AVSS 0.357f $ **FLOATING
C2241 a_23600_43044# AVSS 0.361f $ **FLOATING
C2242 a_19928_43044# AVSS 0.38f $ **FLOATING
C2243 a_18560_43044# AVSS 0.38f $ **FLOATING
C2244 a_14888_43044# AVSS 0.38f $ **FLOATING
C2245 a_13520_43044# AVSS 0.38f $ **FLOATING
C2246 a_9848_43044# AVSS 0.379f $ **FLOATING
C2247 a_8480_43044# AVSS 0.378f $ **FLOATING
C2248 a_4808_43044# AVSS 0.379f $ **FLOATING
C2249 a_3440_43044# AVSS 0.378f $ **FLOATING
C2250 a_n232_43044# AVSS 0.38f $ **FLOATING
C2251 a_23600_43396# AVSS 0.358f $ **FLOATING
C2252 a_19928_43396# AVSS 0.362f $ **FLOATING
C2253 a_18560_43396# AVSS 0.363f $ **FLOATING
C2254 a_14888_43396# AVSS 0.363f $ **FLOATING
C2255 a_13520_43396# AVSS 0.363f $ **FLOATING
C2256 a_9848_43396# AVSS 0.362f $ **FLOATING
C2257 a_8480_43396# AVSS 0.361f $ **FLOATING
C2258 a_4808_43396# AVSS 0.362f $ **FLOATING
C2259 a_3440_43396# AVSS 0.361f $ **FLOATING
C2260 a_n232_43396# AVSS 0.363f $ **FLOATING
C2261 XA8.XA1.XA5.MN0.D AVSS 0.134f
C2262 XA8.XA1.XA2.MN0.D AVSS 1.42f
C2263 XA7.XA1.XA5.MN0.D AVSS 0.15f
C2264 XA7.XA1.XA2.MN0.D AVSS 1.41f
C2265 XA6.XA1.XA5.MN0.D AVSS 0.15f
C2266 XA6.XA1.XA2.MN0.D AVSS 1.41f
C2267 XA5.XA1.XA5.MN0.D AVSS 0.15f
C2268 XA5.XA1.XA2.MN0.D AVSS 1.41f
C2269 XA4.XA1.XA5.MN0.D AVSS 0.15f
C2270 XA4.XA1.XA2.MN0.D AVSS 1.41f
C2271 XA3.XA1.XA5.MN0.D AVSS 0.15f
C2272 XA3.XA1.XA2.MN0.D AVSS 1.41f
C2273 XA2.XA1.XA5.MN0.D AVSS 0.15f
C2274 XA2.XA1.XA2.MN0.D AVSS 1.41f
C2275 XA1.XA1.XA5.MN0.D AVSS 0.15f
C2276 XA1.XA1.XA2.MN0.D AVSS 1.4f
C2277 XA0.XA1.XA5.MN0.D AVSS 0.15f
C2278 XA0.XA1.XA2.MN0.D AVSS 1.41f
C2279 a_23600_43748# AVSS 0.357f $ **FLOATING
C2280 a_19928_43748# AVSS 0.359f $ **FLOATING
C2281 a_18560_43748# AVSS 0.36f $ **FLOATING
C2282 a_14888_43748# AVSS 0.36f $ **FLOATING
C2283 a_13520_43748# AVSS 0.36f $ **FLOATING
C2284 a_9848_43748# AVSS 0.359f $ **FLOATING
C2285 a_8480_43748# AVSS 0.359f $ **FLOATING
C2286 a_4808_43748# AVSS 0.359f $ **FLOATING
C2287 a_3440_43748# AVSS 0.358f $ **FLOATING
C2288 a_n232_43748# AVSS 0.36f $ **FLOATING
C2289 XA8.XA1.XA5.MN1.D AVSS 0.108f
C2290 XA7.XA1.XA5.MN1.D AVSS 0.113f
C2291 XA6.XA1.XA5.MN1.D AVSS 0.113f
C2292 XA5.XA1.XA5.MN1.D AVSS 0.113f
C2293 XA4.XA1.XA5.MN1.D AVSS 0.113f
C2294 XA3.XA1.XA5.MN1.D AVSS 0.113f
C2295 XA2.XA1.XA5.MN1.D AVSS 0.113f
C2296 XA1.XA1.XA5.MN1.D AVSS 0.113f
C2297 XA0.XA1.XA5.MN1.D AVSS 0.113f
C2298 EN AVSS 8.08f
C2299 a_23600_44100# AVSS 0.357f $ **FLOATING
C2300 a_19928_44100# AVSS 0.382f $ **FLOATING
C2301 a_18560_44100# AVSS 0.382f $ **FLOATING
C2302 a_14888_44100# AVSS 0.382f $ **FLOATING
C2303 a_13520_44100# AVSS 0.382f $ **FLOATING
C2304 a_9848_44100# AVSS 0.382f $ **FLOATING
C2305 a_8480_44100# AVSS 0.381f $ **FLOATING
C2306 a_4808_44100# AVSS 0.381f $ **FLOATING
C2307 a_3440_44100# AVSS 0.38f $ **FLOATING
C2308 a_n232_44100# AVSS 0.382f $ **FLOATING
C2309 a_23600_44452# AVSS 0.357f $ **FLOATING
C2310 a_19928_44452# AVSS 0.366f $ **FLOATING
C2311 a_18560_44452# AVSS 0.366f $ **FLOATING
C2312 a_14888_44452# AVSS 0.366f $ **FLOATING
C2313 a_13520_44452# AVSS 0.366f $ **FLOATING
C2314 a_9848_44452# AVSS 0.365f $ **FLOATING
C2315 a_8480_44452# AVSS 0.364f $ **FLOATING
C2316 a_4808_44452# AVSS 0.365f $ **FLOATING
C2317 a_3440_44452# AVSS 0.364f $ **FLOATING
C2318 a_n232_44452# AVSS 0.366f $ **FLOATING
C2319 SARP AVSS 0.301p
C2320 a_23600_44804# AVSS 0.359f $ **FLOATING
C2321 a_19928_44804# AVSS 0.414f $ **FLOATING
C2322 a_18560_44804# AVSS 0.414f $ **FLOATING
C2323 a_14888_44804# AVSS 0.414f $ **FLOATING
C2324 a_13520_44804# AVSS 0.414f $ **FLOATING
C2325 a_9848_44804# AVSS 0.413f $ **FLOATING
C2326 a_8480_44804# AVSS 0.413f $ **FLOATING
C2327 a_4808_44804# AVSS 0.413f $ **FLOATING
C2328 a_3440_44804# AVSS 0.412f $ **FLOATING
C2329 a_n232_44804# AVSS 0.414f $ **FLOATING
C2330 XA20.XA2.MN1.D AVSS 0.573f
C2331 a_23600_45156# AVSS 0.38f $ **FLOATING
C2332 a_19928_45156# AVSS 0.366f $ **FLOATING
C2333 a_18560_45156# AVSS 0.366f $ **FLOATING
C2334 a_14888_45156# AVSS 0.366f $ **FLOATING
C2335 a_13520_45156# AVSS 0.366f $ **FLOATING
C2336 a_9848_45156# AVSS 0.365f $ **FLOATING
C2337 a_8480_45156# AVSS 0.364f $ **FLOATING
C2338 a_4808_45156# AVSS 0.365f $ **FLOATING
C2339 a_3440_45156# AVSS 0.364f $ **FLOATING
C2340 a_n232_45156# AVSS 0.366f $ **FLOATING
C2341 XA8.XA1.XA5.MN2.D AVSS 2.5f
C2342 XA7.XA1.XA5.MN2.D AVSS 2.49f
C2343 XA6.XA1.XA5.MN2.D AVSS 2.49f
C2344 XA5.XA1.XA5.MN2.D AVSS 2.49f
C2345 XA4.XA1.XA5.MN2.D AVSS 2.48f
C2346 XA3.XA1.XA5.MN2.D AVSS 2.47f
C2347 XA2.XA1.XA5.MN2.D AVSS 2.47f
C2348 XA1.XA1.XA5.MN2.D AVSS 2.46f
C2349 XA0.XA1.XA5.MN2.D AVSS 2.48f
C2350 a_23600_45508# AVSS 0.363f $ **FLOATING
C2351 a_19928_45508# AVSS 0.405f $ **FLOATING
C2352 a_18560_45508# AVSS 0.405f $ **FLOATING
C2353 a_14888_45508# AVSS 0.405f $ **FLOATING
C2354 a_13520_45508# AVSS 0.405f $ **FLOATING
C2355 a_9848_45508# AVSS 0.405f $ **FLOATING
C2356 a_8480_45508# AVSS 0.404f $ **FLOATING
C2357 a_4808_45508# AVSS 0.404f $ **FLOATING
C2358 a_3440_45508# AVSS 0.403f $ **FLOATING
C2359 a_n232_45508# AVSS 0.405f $ **FLOATING
C2360 a_23600_45860# AVSS 0.404f $ **FLOATING
C2361 a_19928_45860# AVSS 0.366f $ **FLOATING
C2362 a_18560_45860# AVSS 0.366f $ **FLOATING
C2363 a_14888_45860# AVSS 0.366f $ **FLOATING
C2364 a_13520_45860# AVSS 0.366f $ **FLOATING
C2365 a_9848_45860# AVSS 0.366f $ **FLOATING
C2366 a_8480_45860# AVSS 0.366f $ **FLOATING
C2367 a_4808_45860# AVSS 0.366f $ **FLOATING
C2368 a_3440_45860# AVSS 0.366f $ **FLOATING
C2369 a_n232_45860# AVSS 0.366f $ **FLOATING
C2370 a_23600_46212# AVSS 0.368f $ **FLOATING
C2371 a_19928_46212# AVSS 0.415f $ **FLOATING
C2372 a_18560_46212# AVSS 0.415f $ **FLOATING
C2373 a_14888_46212# AVSS 0.415f $ **FLOATING
C2374 a_13520_46212# AVSS 0.415f $ **FLOATING
C2375 a_9848_46212# AVSS 0.415f $ **FLOATING
C2376 a_8480_46212# AVSS 0.415f $ **FLOATING
C2377 a_4808_46212# AVSS 0.415f $ **FLOATING
C2378 a_3440_46212# AVSS 0.415f $ **FLOATING
C2379 a_n232_46212# AVSS 0.416f $ **FLOATING
C2380 XA20.XA2a.MN0.D AVSS 17.9f
C2381 a_23600_46564# AVSS 0.404f $ **FLOATING
C2382 a_19928_46564# AVSS 0.366f $ **FLOATING
C2383 a_18560_46564# AVSS 0.366f $ **FLOATING
C2384 a_14888_46564# AVSS 0.366f $ **FLOATING
C2385 a_13520_46564# AVSS 0.366f $ **FLOATING
C2386 a_9848_46564# AVSS 0.366f $ **FLOATING
C2387 a_8480_46564# AVSS 0.366f $ **FLOATING
C2388 a_4808_46564# AVSS 0.366f $ **FLOATING
C2389 a_3440_46564# AVSS 0.366f $ **FLOATING
C2390 a_n232_46564# AVSS 0.366f $ **FLOATING
C2391 XA8.XA3.MN0.G AVSS 3.68f
C2392 XA7.XA3.MN0.G AVSS 3.66f
C2393 XA6.XA3.MN0.G AVSS 3.66f
C2394 XA5.XA3.MN0.G AVSS 3.66f
C2395 XA4.XA3.MN0.G AVSS 3.66f
C2396 XA3.XA3.MN0.G AVSS 11f
C2397 XA2.XA3.MN0.G AVSS 11.1f
C2398 XA1.XA3.MN0.G AVSS 10.4f
C2399 D<8> AVSS 19.5f
C2400 a_23600_46916# AVSS 0.368f $ **FLOATING
C2401 a_19928_46916# AVSS 0.406f $ **FLOATING
C2402 a_18560_46916# AVSS 0.406f $ **FLOATING
C2403 a_14888_46916# AVSS 0.406f $ **FLOATING
C2404 a_13520_46916# AVSS 0.406f $ **FLOATING
C2405 a_9848_46916# AVSS 0.406f $ **FLOATING
C2406 a_8480_46916# AVSS 0.406f $ **FLOATING
C2407 a_4808_46916# AVSS 0.406f $ **FLOATING
C2408 a_3440_46916# AVSS 0.406f $ **FLOATING
C2409 a_n232_46916# AVSS 0.406f $ **FLOATING
C2410 a_23600_47268# AVSS 0.404f $ **FLOATING
C2411 a_19928_47268# AVSS 0.366f $ **FLOATING
C2412 a_18560_47268# AVSS 0.366f $ **FLOATING
C2413 a_14888_47268# AVSS 0.366f $ **FLOATING
C2414 a_13520_47268# AVSS 0.366f $ **FLOATING
C2415 a_9848_47268# AVSS 0.366f $ **FLOATING
C2416 a_8480_47268# AVSS 0.366f $ **FLOATING
C2417 a_4808_47268# AVSS 0.366f $ **FLOATING
C2418 a_3440_47268# AVSS 0.366f $ **FLOATING
C2419 a_n232_47268# AVSS 0.366f $ **FLOATING
C2420 a_23600_47620# AVSS 0.368f $ **FLOATING
C2421 a_19928_47620# AVSS 0.414f $ **FLOATING
C2422 a_18560_47620# AVSS 0.414f $ **FLOATING
C2423 a_14888_47620# AVSS 0.414f $ **FLOATING
C2424 a_13520_47620# AVSS 0.414f $ **FLOATING
C2425 a_9848_47620# AVSS 0.414f $ **FLOATING
C2426 a_8480_47620# AVSS 0.414f $ **FLOATING
C2427 a_4808_47620# AVSS 0.414f $ **FLOATING
C2428 a_3440_47620# AVSS 0.414f $ **FLOATING
C2429 a_n232_47620# AVSS 0.414f $ **FLOATING
C2430 XA20.XA3a.MN0.D AVSS 22.7f
C2431 a_23600_47972# AVSS 0.404f $ **FLOATING
C2432 a_19928_47972# AVSS 0.366f $ **FLOATING
C2433 a_18560_47972# AVSS 0.366f $ **FLOATING
C2434 a_14888_47972# AVSS 0.366f $ **FLOATING
C2435 a_13520_47972# AVSS 0.366f $ **FLOATING
C2436 a_9848_47972# AVSS 0.366f $ **FLOATING
C2437 a_8480_47972# AVSS 0.366f $ **FLOATING
C2438 a_4808_47972# AVSS 0.366f $ **FLOATING
C2439 a_3440_47972# AVSS 0.366f $ **FLOATING
C2440 a_n232_47972# AVSS 0.366f $ **FLOATING
C2441 XA8.XA4.MN0.G AVSS 3.84f
C2442 XA7.XA4.MN0.G AVSS 3.82f
C2443 XA6.XA4.MN0.G AVSS 3.82f
C2444 XA5.XA4.MN0.G AVSS 3.82f
C2445 XA4.XA4.MN0.G AVSS 3.82f
C2446 XA3.XA4.MN0.G AVSS 3.81f
C2447 XA2.XA4.MN0.G AVSS 3.82f
C2448 XA1.XA4.MN0.G AVSS 3.81f
C2449 XA0.XA4.MN0.G AVSS 3.96f
C2450 a_23600_48324# AVSS 0.362f $ **FLOATING
C2451 a_19928_48324# AVSS 0.405f $ **FLOATING
C2452 a_18560_48324# AVSS 0.405f $ **FLOATING
C2453 a_14888_48324# AVSS 0.405f $ **FLOATING
C2454 a_13520_48324# AVSS 0.405f $ **FLOATING
C2455 a_9848_48324# AVSS 0.405f $ **FLOATING
C2456 a_8480_48324# AVSS 0.405f $ **FLOATING
C2457 a_4808_48324# AVSS 0.405f $ **FLOATING
C2458 a_3440_48324# AVSS 0.405f $ **FLOATING
C2459 a_n232_48324# AVSS 0.405f $ **FLOATING
C2460 a_23600_48676# AVSS 0.358f $ **FLOATING
C2461 a_19928_48676# AVSS 0.366f $ **FLOATING
C2462 a_18560_48676# AVSS 0.366f $ **FLOATING
C2463 a_14888_48676# AVSS 0.366f $ **FLOATING
C2464 a_13520_48676# AVSS 0.366f $ **FLOATING
C2465 a_9848_48676# AVSS 0.366f $ **FLOATING
C2466 a_8480_48676# AVSS 0.366f $ **FLOATING
C2467 a_4808_48676# AVSS 0.366f $ **FLOATING
C2468 a_3440_48676# AVSS 0.366f $ **FLOATING
C2469 a_n232_48676# AVSS 0.366f $ **FLOATING
C2470 a_23600_49028# AVSS 0.357f $ **FLOATING
C2471 a_19928_49028# AVSS 0.416f $ **FLOATING
C2472 a_18560_49028# AVSS 0.416f $ **FLOATING
C2473 a_14888_49028# AVSS 0.416f $ **FLOATING
C2474 a_13520_49028# AVSS 0.416f $ **FLOATING
C2475 a_9848_49028# AVSS 0.416f $ **FLOATING
C2476 a_8480_49028# AVSS 0.416f $ **FLOATING
C2477 a_4808_49028# AVSS 0.416f $ **FLOATING
C2478 a_3440_49028# AVSS 0.416f $ **FLOATING
C2479 a_n232_49028# AVSS 0.416f $ **FLOATING
C2480 a_23600_49380# AVSS 0.357f $ **FLOATING
C2481 a_19928_49380# AVSS 0.366f $ **FLOATING
C2482 a_18560_49380# AVSS 0.366f $ **FLOATING
C2483 a_14888_49380# AVSS 0.366f $ **FLOATING
C2484 a_13520_49380# AVSS 0.366f $ **FLOATING
C2485 a_9848_49380# AVSS 0.366f $ **FLOATING
C2486 a_8480_49380# AVSS 0.366f $ **FLOATING
C2487 a_4808_49380# AVSS 0.366f $ **FLOATING
C2488 a_3440_49380# AVSS 0.366f $ **FLOATING
C2489 a_n232_49380# AVSS 0.366f $ **FLOATING
C2490 XA8.XA4.MN0.D AVSS 3.72f
C2491 XA7.XA4.MN0.D AVSS 3.72f
C2492 XA6.XA4.MN0.D AVSS 3.72f
C2493 XA5.XA4.MN0.D AVSS 3.72f
C2494 XA4.XA4.MN0.D AVSS 3.72f
C2495 XA3.XA4.MN0.D AVSS 6.94f
C2496 XA2.XA4.MN0.D AVSS 7.16f
C2497 XA1.XA4.MN0.D AVSS 12.6f
C2498 VREF AVSS 27.8f
C2499 XA0.XA4.MN0.D AVSS 17.4f
C2500 a_23600_49732# AVSS 0.358f $ **FLOATING
C2501 a_19928_49732# AVSS 0.406f $ **FLOATING
C2502 a_18560_49732# AVSS 0.406f $ **FLOATING
C2503 a_14888_49732# AVSS 0.406f $ **FLOATING
C2504 a_13520_49732# AVSS 0.406f $ **FLOATING
C2505 a_9848_49732# AVSS 0.406f $ **FLOATING
C2506 a_8480_49732# AVSS 0.406f $ **FLOATING
C2507 a_4808_49732# AVSS 0.406f $ **FLOATING
C2508 a_3440_49732# AVSS 0.406f $ **FLOATING
C2509 a_n232_49732# AVSS 0.406f $ **FLOATING
C2510 XA20.XA3.MN0.D AVSS 2.31f
C2511 a_23600_50084# AVSS 0.359f $ **FLOATING
C2512 a_19928_50084# AVSS 0.366f $ **FLOATING
C2513 a_18560_50084# AVSS 0.363f $ **FLOATING
C2514 a_14888_50084# AVSS 0.363f $ **FLOATING
C2515 a_13520_50084# AVSS 0.363f $ **FLOATING
C2516 a_9848_50084# AVSS 0.363f $ **FLOATING
C2517 a_8480_50084# AVSS 0.363f $ **FLOATING
C2518 a_4808_50084# AVSS 0.363f $ **FLOATING
C2519 a_3440_50084# AVSS 0.363f $ **FLOATING
C2520 a_n232_50084# AVSS 0.363f $ **FLOATING
C2521 XA20.XA3.MN1.D AVSS 0.597f
C2522 XA20.XA3.MN6.D AVSS 3.02f
C2523 XA20.XA3a.MN0.G AVSS 2.98f
C2524 XA8.XA6.MN0.D AVSS 0.218f
C2525 XA8.XA6.MP0.G AVSS 0.964f
C2526 XA7.XA6.MN0.D AVSS 0.201f
C2527 XA7.XA6.MP0.G AVSS 8.77f
C2528 XA6.XA6.MN0.D AVSS 0.201f
C2529 XA6.XA6.MP0.G AVSS 6.39f
C2530 XA5.XA6.MN0.D AVSS 0.201f
C2531 XA5.XA6.MP0.G AVSS 5.21f
C2532 XA4.XA6.MN0.D AVSS 0.201f
C2533 XA4.XA6.MP0.G AVSS 6.53f
C2534 XA3.XA6.MN0.D AVSS 0.201f
C2535 XA3.XA6.MP0.G AVSS 4.62f
C2536 XA2.XA6.MN0.D AVSS 0.201f
C2537 XA2.XA6.MP0.G AVSS 4.95f
C2538 XA1.XA6.MN0.D AVSS 0.201f
C2539 XA1.XA6.MP0.G AVSS 10.6f
C2540 XA0.XA6.MN0.D AVSS 0.201f
C2541 XA0.XA6.MP0.G AVSS 15.1f
C2542 a_23600_50436# AVSS 0.381f $ **FLOATING
C2543 a_19928_50436# AVSS 0.416f $ **FLOATING
C2544 a_18560_50436# AVSS 0.415f $ **FLOATING
C2545 a_14888_50436# AVSS 0.415f $ **FLOATING
C2546 a_13520_50436# AVSS 0.415f $ **FLOATING
C2547 a_9848_50436# AVSS 0.415f $ **FLOATING
C2548 a_8480_50436# AVSS 0.415f $ **FLOATING
C2549 a_4808_50436# AVSS 0.415f $ **FLOATING
C2550 a_3440_50436# AVSS 0.415f $ **FLOATING
C2551 a_n232_50436# AVSS 0.416f $ **FLOATING
C2552 a_23600_50788# AVSS 0.361f $ **FLOATING
C2553 a_19928_50788# AVSS 0.361f $ **FLOATING
C2554 a_18560_50788# AVSS 0.363f $ **FLOATING
C2555 a_14888_50788# AVSS 0.363f $ **FLOATING
C2556 a_13520_50788# AVSS 0.363f $ **FLOATING
C2557 a_9848_50788# AVSS 0.363f $ **FLOATING
C2558 a_8480_50788# AVSS 0.363f $ **FLOATING
C2559 a_4808_50788# AVSS 0.363f $ **FLOATING
C2560 a_3440_50788# AVSS 0.363f $ **FLOATING
C2561 a_n232_50788# AVSS 0.363f $ **FLOATING
C2562 XA8.XA6.MN2.D AVSS 0.141f
C2563 D<0> AVSS 1.24f
C2564 XA7.XA6.MN2.D AVSS 0.15f
C2565 D<1> AVSS 11.9f
C2566 XA6.XA6.MN2.D AVSS 0.15f
C2567 D<2> AVSS 9.38f
C2568 XA5.XA6.MN2.D AVSS 0.15f
C2569 D<3> AVSS 8.3f
C2570 XA4.XA6.MN2.D AVSS 0.15f
C2571 D<4> AVSS 8.94f
C2572 XA3.XA6.MN2.D AVSS 0.15f
C2573 D<5> AVSS 8.41f
C2574 XA2.XA6.MN2.D AVSS 0.15f
C2575 D<6> AVSS 9.43f
C2576 XA1.XA6.MN2.D AVSS 0.15f
C2577 D<7> AVSS 8.44f
C2578 XA0.XA6.MN2.D AVSS 0.15f
C2579 XA0.XA6.MP2.G AVSS 14.9f
C2580 a_23600_51140# AVSS 0.358f $ **FLOATING
C2581 a_19928_51140# AVSS 0.382f $ **FLOATING
C2582 a_18560_51140# AVSS 0.383f $ **FLOATING
C2583 a_14888_51140# AVSS 0.383f $ **FLOATING
C2584 a_13520_51140# AVSS 0.383f $ **FLOATING
C2585 a_9848_51140# AVSS 0.383f $ **FLOATING
C2586 a_8480_51140# AVSS 0.383f $ **FLOATING
C2587 a_4808_51140# AVSS 0.383f $ **FLOATING
C2588 a_3440_51140# AVSS 0.383f $ **FLOATING
C2589 a_n232_51140# AVSS 0.383f $ **FLOATING
C2590 XA8.XA7.MN0.G AVSS 1.85f
C2591 XA8.XA1.XA5.MN2.G AVSS 4.7f
C2592 XA7.XA1.XA5.MN2.G AVSS 4.58f
C2593 XA6.XA1.XA5.MN2.G AVSS 4.65f
C2594 XA5.XA1.XA5.MN2.G AVSS 4.59f
C2595 XA4.XA1.XA5.MN2.G AVSS 4.67f
C2596 XA3.XA1.XA5.MN2.G AVSS 4.64f
C2597 XA2.XA1.XA5.MN2.G AVSS 4.63f
C2598 XA0.XA7.MN0.G AVSS 4.64f
C2599 a_23600_51492# AVSS 0.357f $ **FLOATING
C2600 a_19928_51492# AVSS 0.387f $ **FLOATING
C2601 a_18560_51492# AVSS 0.387f $ **FLOATING
C2602 a_14888_51492# AVSS 0.387f $ **FLOATING
C2603 a_13520_51492# AVSS 0.387f $ **FLOATING
C2604 a_9848_51492# AVSS 0.387f $ **FLOATING
C2605 a_8480_51492# AVSS 0.387f $ **FLOATING
C2606 a_4808_51492# AVSS 0.387f $ **FLOATING
C2607 a_3440_51492# AVSS 0.387f $ **FLOATING
C2608 a_n232_51492# AVSS 0.388f $ **FLOATING
C2609 XA7.XA8.MN0.D AVSS 0.223f
C2610 XA6.XA8.MN0.D AVSS 0.223f
C2611 XA5.XA8.MN0.D AVSS 0.223f
C2612 XA4.XA8.MN0.D AVSS 0.223f
C2613 XA3.XA8.MN0.D AVSS 0.223f
C2614 XA2.XA8.MN0.D AVSS 0.223f
C2615 XA1.XA8.MN0.D AVSS 0.223f
C2616 XA0.XA8.MN0.D AVSS 0.223f
C2617 a_23600_51844# AVSS 0.357f $ **FLOATING
C2618 a_19928_51844# AVSS 0.384f $ **FLOATING
C2619 a_18560_51844# AVSS 0.386f $ **FLOATING
C2620 a_14888_51844# AVSS 0.386f $ **FLOATING
C2621 a_13520_51844# AVSS 0.386f $ **FLOATING
C2622 a_9848_51844# AVSS 0.386f $ **FLOATING
C2623 a_8480_51844# AVSS 0.386f $ **FLOATING
C2624 a_4808_51844# AVSS 0.386f $ **FLOATING
C2625 a_3440_51844# AVSS 0.386f $ **FLOATING
C2626 a_n232_51844# AVSS 0.386f $ **FLOATING
C2627 XA8.XA7.MN0.D AVSS 1.52f
C2628 XA7.XA7.MN0.D AVSS 1.53f
C2629 XA6.XA7.MN0.D AVSS 1.53f
C2630 XA5.XA7.MN0.D AVSS 1.53f
C2631 XA4.XA7.MN0.D AVSS 1.53f
C2632 XA3.XA7.MN0.D AVSS 1.53f
C2633 XA2.XA7.MN0.D AVSS 1.53f
C2634 XA1.XA7.MN0.D AVSS 1.53f
C2635 XA0.XA7.MN0.D AVSS 1.53f
C2636 a_23600_52196# AVSS 0.357f $ **FLOATING
C2637 a_19928_52196# AVSS 0.364f $ **FLOATING
C2638 a_18560_52196# AVSS 0.364f $ **FLOATING
C2639 a_14888_52196# AVSS 0.364f $ **FLOATING
C2640 a_13520_52196# AVSS 0.364f $ **FLOATING
C2641 a_9848_52196# AVSS 0.364f $ **FLOATING
C2642 a_8480_52196# AVSS 0.364f $ **FLOATING
C2643 a_4808_52196# AVSS 0.364f $ **FLOATING
C2644 a_3440_52196# AVSS 0.364f $ **FLOATING
C2645 a_n232_52196# AVSS 0.365f $ **FLOATING
C2646 SARN AVSS 0.302p
C2647 XA8.XA9.MN0.D AVSS 0.174f
C2648 XA8.XA9.MN1.G AVSS 1.72f
C2649 XA7.XA9.MN0.D AVSS 0.174f
C2650 XA7.XA9.MN1.G AVSS 1.73f
C2651 XA6.XA9.MN0.D AVSS 0.174f
C2652 XA6.XA9.MN1.G AVSS 1.74f
C2653 XA5.XA9.MN0.D AVSS 0.174f
C2654 XA5.XA9.MN1.G AVSS 1.73f
C2655 XA4.XA9.MN0.D AVSS 0.174f
C2656 XA4.XA9.MN1.G AVSS 1.74f
C2657 XA3.XA9.MN0.D AVSS 0.174f
C2658 XA3.XA9.MN1.G AVSS 1.73f
C2659 XA2.XA9.MN0.D AVSS 0.174f
C2660 XA2.XA9.MN1.G AVSS 1.74f
C2661 XA1.XA9.MN0.D AVSS 0.174f
C2662 XA1.XA9.MN1.G AVSS 1.73f
C2663 XA0.XA9.MN0.D AVSS 0.174f
C2664 XA0.XA9.MN1.G AVSS 1.8f
C2665 a_23600_52548# AVSS 0.359f $ **FLOATING
C2666 a_19928_52548# AVSS 0.383f $ **FLOATING
C2667 a_18560_52548# AVSS 0.383f $ **FLOATING
C2668 a_14888_52548# AVSS 0.383f $ **FLOATING
C2669 a_13520_52548# AVSS 0.383f $ **FLOATING
C2670 a_9848_52548# AVSS 0.383f $ **FLOATING
C2671 a_8480_52548# AVSS 0.383f $ **FLOATING
C2672 a_4808_52548# AVSS 0.383f $ **FLOATING
C2673 a_3440_52548# AVSS 0.383f $ **FLOATING
C2674 a_n232_52548# AVSS 0.383f $ **FLOATING
C2675 XA20.XA4.MN0.D AVSS 0.862f
C2676 XA8.XA10.MN0.G AVSS 0.929f
C2677 XA7.XA10.MN0.G AVSS 0.929f
C2678 XA6.XA10.MN0.G AVSS 0.929f
C2679 XA5.XA10.MN0.G AVSS 0.929f
C2680 XA4.XA10.MN0.G AVSS 0.929f
C2681 XA3.XA10.MN0.G AVSS 0.929f
C2682 XA2.XA10.MN0.G AVSS 0.929f
C2683 XA1.XA10.MN0.G AVSS 0.929f
C2684 XA0.XA10.MN0.G AVSS 0.929f
C2685 a_23600_52900# AVSS 0.382f $ **FLOATING
C2686 a_19928_52900# AVSS 0.387f $ **FLOATING
C2687 a_18560_52900# AVSS 0.387f $ **FLOATING
C2688 a_14888_52900# AVSS 0.387f $ **FLOATING
C2689 a_13520_52900# AVSS 0.387f $ **FLOATING
C2690 a_9848_52900# AVSS 0.387f $ **FLOATING
C2691 a_8480_52900# AVSS 0.387f $ **FLOATING
C2692 a_4808_52900# AVSS 0.387f $ **FLOATING
C2693 a_3440_52900# AVSS 0.387f $ **FLOATING
C2694 a_n232_52900# AVSS 0.388f $ **FLOATING
C2695 XA20.XA9.MN0.D AVSS 6.27f
C2696 XA8.XA10.MN0.D AVSS 0.902f
C2697 XA7.XA10.MN0.D AVSS 0.9f
C2698 XA6.XA10.MN0.D AVSS 0.902f
C2699 XA5.XA10.MN0.D AVSS 0.9f
C2700 XA4.XA10.MN0.D AVSS 0.902f
C2701 XA3.XA10.MN0.D AVSS 0.9f
C2702 XA2.XA10.MN0.D AVSS 0.902f
C2703 XA1.XA10.MN0.D AVSS 0.9f
C2704 XA0.XA10.MN0.D AVSS 0.902f
C2705 a_23600_53252# AVSS 0.388f $ **FLOATING
C2706 a_19928_53252# AVSS 0.371f $ **FLOATING
C2707 a_18560_53252# AVSS 0.365f $ **FLOATING
C2708 a_14888_53252# AVSS 0.371f $ **FLOATING
C2709 a_13520_53252# AVSS 0.365f $ **FLOATING
C2710 a_9848_53252# AVSS 0.371f $ **FLOATING
C2711 a_8480_53252# AVSS 0.365f $ **FLOATING
C2712 a_4808_53252# AVSS 0.371f $ **FLOATING
C2713 a_3440_53252# AVSS 0.365f $ **FLOATING
C2714 a_n232_53252# AVSS 0.371f $ **FLOATING
C2715 XA0.XA11.MN1.G AVSS 42.4f
C2716 a_23600_53604# AVSS 0.363f $ **FLOATING
C2717 a_19928_53604# AVSS 0.406f $ **FLOATING
C2718 a_18560_53604# AVSS 0.405f $ **FLOATING
C2719 a_14888_53604# AVSS 0.406f $ **FLOATING
C2720 a_13520_53604# AVSS 0.405f $ **FLOATING
C2721 a_9848_53604# AVSS 0.406f $ **FLOATING
C2722 a_8480_53604# AVSS 0.405f $ **FLOATING
C2723 a_4808_53604# AVSS 0.406f $ **FLOATING
C2724 a_3440_53604# AVSS 0.405f $ **FLOATING
C2725 a_n232_53604# AVSS 0.406f $ **FLOATING
C2726 XA20.XA10.MN0.D AVSS 0.136f
C2727 XA20.XA10.MN1.D AVSS 7.1f
C2728 XA8.XA12.MN0.G AVSS 1.18f
C2729 XA7.XA12.MN0.G AVSS 1.14f
C2730 XA8.XA11.MN1.G AVSS 1.7f
C2731 XA6.XA12.MN0.G AVSS 1.18f
C2732 XA7.XA11.MN1.G AVSS 1.55f
C2733 XA5.XA12.MN0.G AVSS 1.14f
C2734 XA6.XA11.MN1.G AVSS 1.7f
C2735 XA4.XA12.MN0.G AVSS 1.18f
C2736 XA5.XA11.MN1.G AVSS 1.55f
C2737 XA3.XA12.MN0.G AVSS 1.14f
C2738 XA4.XA11.MN1.G AVSS 1.7f
C2739 XA2.XA12.MN0.G AVSS 1.18f
C2740 XA3.XA11.MN1.G AVSS 1.55f
C2741 XA1.XA12.MN0.G AVSS 1.14f
C2742 XA2.XA11.MN1.G AVSS 1.7f
C2743 XA0.XA12.MN0.G AVSS 1.18f
C2744 XA0.XA12.MN0.D AVSS 1.55f
C2745 a_23600_53956# AVSS 0.383f $ **FLOATING
C2746 a_19928_53956# AVSS 0.47f $ **FLOATING
C2747 a_18560_53956# AVSS 0.471f $ **FLOATING
C2748 a_14888_53956# AVSS 0.47f $ **FLOATING
C2749 a_13520_53956# AVSS 0.471f $ **FLOATING
C2750 a_9848_53956# AVSS 0.47f $ **FLOATING
C2751 a_8480_53956# AVSS 0.471f $ **FLOATING
C2752 a_4808_53956# AVSS 0.47f $ **FLOATING
C2753 a_3440_53956# AVSS 0.471f $ **FLOATING
C2754 a_n232_53956# AVSS 0.47f $ **FLOATING
C2755 CK_SAMPLE AVSS 23.5f
C2756 a_23600_54308# AVSS 0.37f $ **FLOATING
C2757 a_19928_54308# AVSS 0.539f $ **FLOATING
C2758 a_18560_54308# AVSS 0.538f $ **FLOATING
C2759 a_14888_54308# AVSS 0.539f $ **FLOATING
C2760 a_13520_54308# AVSS 0.538f $ **FLOATING
C2761 a_9848_54308# AVSS 0.539f $ **FLOATING
C2762 a_8480_54308# AVSS 0.538f $ **FLOATING
C2763 a_4808_54308# AVSS 0.539f $ **FLOATING
C2764 a_3440_54308# AVSS 0.538f $ **FLOATING
C2765 a_n232_54308# AVSS 0.539f $ **FLOATING
C2766 DONE AVSS 1.18f
C2767 XA20.XA11.MN0.D AVSS 1.24f
C2768 a_23600_54660# AVSS 0.407f $ **FLOATING
C2769 XA20.XA12.MN0.G AVSS 1.12f
C2770 XA20.XA12.MN0.D AVSS 0.791f
C2771 a_23600_55012# AVSS 0.471f $ **FLOATING
C2772 a_23600_55364# AVSS 0.541f $ **FLOATING
C2773 AVDD AVSS 0.691p
.ends

