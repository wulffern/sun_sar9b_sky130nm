magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 1260 4928
<< locali >>
rect 828 1435 912 1469
rect 912 2887 1044 2921
rect 912 2095 1044 2129
rect 912 1435 946 2921
rect 98 775 216 809
rect 98 951 216 985
rect 98 2535 216 2569
rect 98 3767 216 3801
rect 98 775 132 3801
rect 216 3767 300 3801
rect 300 3987 432 4021
rect 300 3767 334 4021
rect 314 4427 432 4461
rect 216 4119 314 4153
rect 314 4119 348 4461
rect 828 4691 912 4725
rect 912 4207 1044 4241
rect 912 4207 946 4725
rect 314 1347 432 1381
rect 314 2931 432 2965
rect 314 1347 348 2965
rect 162 4383 270 4417
rect 162 4647 270 4681
rect 162 4471 270 4505
rect 378 2139 486 2173
rect 378 1699 486 1733
rect 162 687 270 721
rect 162 2975 270 3009
<< m1 >>
rect 828 2843 912 2877
rect 912 1391 1044 1425
rect 912 1655 1044 1689
rect 912 1391 946 2877
rect 216 687 300 721
rect 216 1039 300 1073
rect 300 687 334 1073
rect 216 2975 300 3009
rect 216 3327 300 3361
rect 300 2975 334 3361
rect 98 247 216 281
rect 98 3239 216 3273
rect 98 3943 216 3977
rect 98 247 132 3977
rect 216 3943 300 3977
rect 300 4251 432 4285
rect 300 3943 334 4285
<< m3 >>
rect 774 0 866 4928
rect 378 0 470 4928
rect 774 0 866 4928
rect 378 0 470 4928
use SUNSAR_TAPCELLB_CV XA0 
transform 1 0 0 0 1 0
box 0 0 1260 176
use SUNSAR_SARKICKHX1_CV XA1 
transform 1 0 0 0 1 176
box 0 176 1260 880
use SUNSAR_SARCMPHX1_CV XA2 
transform 1 0 0 0 1 880
box 0 880 1260 1584
use SUNSAR_IVX4_CV XA2a 
transform 1 0 0 0 1 1584
box 0 1584 1260 2024
use SUNSAR_IVX4_CV XA3a 
transform 1 0 0 0 1 2024
box 0 2024 1260 2464
use SUNSAR_SARCMPHX1_CV XA3 
transform 1 0 0 0 1 2464
box 0 2464 1260 3168
use SUNSAR_SARKICKHX1_CV XA4 
transform 1 0 0 0 1 3168
box 0 3168 1260 3872
use SUNSAR_IVX1_CV XA9 
transform 1 0 0 0 1 3872
box 0 3872 1260 4048
use SUNSAR_NDX1_CV XA10 
transform 1 0 0 0 1 4048
box 0 4048 1260 4312
use SUNSAR_NRX1_CV XA11 
transform 1 0 0 0 1 4312
box 0 4312 1260 4576
use SUNSAR_IVX1_CV XA12 
transform 1 0 0 0 1 4576
box 0 4576 1260 4752
use SUNSAR_TAPCELLB_CV XA13 
transform 1 0 0 0 1 4752
box 0 4752 1260 4928
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 774 0 1 2843
box 774 2843 866 2877
use SUNSAR_cut_M1M2_2x1 xcut1 
transform 1 0 990 0 1 1391
box 990 1391 1082 1425
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 990 0 1 1655
box 990 1655 1082 1689
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 178 0 1 687
box 178 687 270 721
use SUNSAR_cut_M1M2_2x1 xcut4 
transform 1 0 178 0 1 1039
box 178 1039 270 1073
use SUNSAR_cut_M1M2_2x1 xcut5 
transform 1 0 178 0 1 2975
box 178 2975 270 3009
use SUNSAR_cut_M1M2_2x1 xcut6 
transform 1 0 178 0 1 3327
box 178 3327 270 3361
use SUNSAR_cut_M1M2_2x1 xcut7 
transform 1 0 162 0 1 247
box 162 247 254 281
use SUNSAR_cut_M1M2_2x1 xcut8 
transform 1 0 162 0 1 3239
box 162 3239 254 3273
use SUNSAR_cut_M1M2_2x1 xcut9 
transform 1 0 162 0 1 3943
box 162 3943 254 3977
use SUNSAR_cut_M1M2_2x1 xcut10 
transform 1 0 162 0 1 3943
box 162 3943 254 3977
use SUNSAR_cut_M1M2_2x1 xcut11 
transform 1 0 378 0 1 4251
box 378 4251 470 4285
<< labels >>
flabel locali s 162 4383 270 4417 0 FreeSans 400 0 0 0 CK_SAMPLE
port 6 nsew signal bidirectional
flabel locali s 162 4647 270 4681 0 FreeSans 400 0 0 0 CK_CMP
port 5 nsew signal bidirectional
flabel locali s 162 4471 270 4505 0 FreeSans 400 0 0 0 DONE
port 7 nsew signal bidirectional
flabel locali s 378 2139 486 2173 0 FreeSans 400 0 0 0 CNO
port 4 nsew signal bidirectional
flabel locali s 378 1699 486 1733 0 FreeSans 400 0 0 0 CPO
port 3 nsew signal bidirectional
flabel locali s 162 687 270 721 0 FreeSans 400 0 0 0 CPI
port 1 nsew signal bidirectional
flabel locali s 162 2975 270 3009 0 FreeSans 400 0 0 0 CNI
port 2 nsew signal bidirectional
flabel m3 s 774 0 866 4928 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 378 0 470 4928 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 4928
<< end >>
