magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect 0 0 2520 4224
<< locali >>
rect 2088 498 2256 558
rect 2088 2962 2256 3022
rect 2088 4018 2256 4078
rect 2256 498 2316 4078
rect 480 1846 600 1906
rect 600 1642 864 1702
rect 600 1642 660 1906
rect 480 1906 540 1966
rect 432 3666 600 3726
rect 600 1994 864 2054
rect 600 1994 660 3726
rect 432 2610 600 2670
rect 600 1994 864 2054
rect 600 1994 660 2670
rect 204 850 432 910
rect 204 3314 432 3374
rect 204 850 264 3374
rect 324 2258 540 2318
rect 1980 4018 2196 4078
rect 324 498 540 558
rect 324 3314 540 3374
rect 756 3050 972 3110
rect 756 4106 972 4166
rect 1548 762 1764 822
<< m1 >>
rect 432 1202 600 1262
rect 432 2258 600 2318
rect 600 1202 660 2318
rect 204 498 432 558
rect 204 4018 432 4078
rect 204 2962 432 3022
rect 204 498 264 4078
<< m3 >>
rect 1548 0 1748 4224
rect 756 0 956 4224
rect 1548 0 1748 4224
rect 756 0 956 4224
use SUNSAR_TAPCELLB_CV XA0 
transform 1 0 0 0 1 0
box 0 0 2520 352
use SUNSAR_SAREMX1_CV XA1 
transform 1 0 0 0 1 352
box 0 352 2520 1760
use SUNSAR_IVX1_CV XA2 
transform 1 0 0 0 1 1760
box 0 1760 2520 2112
use SUNSAR_SARLTX1_CV XA4 
transform 1 0 0 0 1 2112
box 0 2112 2520 3168
use SUNSAR_SARLTX1_CV XA5 
transform 1 0 0 0 1 3168
box 0 3168 2520 4224
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 356 0 1 1202
box 356 1202 540 1270
use SUNSAR_cut_M1M2_2x1 xcut1 
transform 1 0 356 0 1 2258
box 356 2258 540 2326
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 324 0 1 498
box 324 498 508 566
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 324 0 1 4018
box 324 4018 508 4086
use SUNSAR_cut_M1M2_2x1 xcut4 
transform 1 0 324 0 1 2962
box 324 2962 508 3030
<< labels >>
flabel locali s 324 2258 540 2318 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew signal bidirectional
flabel locali s 1980 4018 2196 4078 0 FreeSans 400 0 0 0 RST_N
port 4 nsew signal bidirectional
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 EN
port 3 nsew signal bidirectional
flabel locali s 324 3314 540 3374 0 FreeSans 400 0 0 0 CMP_ON
port 2 nsew signal bidirectional
flabel locali s 756 3050 972 3110 0 FreeSans 400 0 0 0 CHL_OP
port 6 nsew signal bidirectional
flabel locali s 756 4106 972 4166 0 FreeSans 400 0 0 0 CHL_ON
port 7 nsew signal bidirectional
flabel locali s 1548 762 1764 822 0 FreeSans 400 0 0 0 ENO
port 5 nsew signal bidirectional
flabel m3 s 1548 0 1748 4224 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 756 0 956 4224 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 2520 0 4224
<< end >>
