magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect 0 0 7272 1056
<< m1 >>
rect 108 -44 7236 44
rect 7164 44 7236 132
rect 108 132 7092 220
rect 7164 132 7236 220
rect 108 220 180 308
rect 7164 220 7236 308
rect 108 308 180 396
rect 252 308 7236 396
rect 108 396 180 484
rect 7164 396 7236 484
rect 108 484 7092 572
rect 7164 484 7236 572
rect 108 572 180 660
rect 7164 572 7236 660
rect 108 660 180 748
rect 252 660 7236 748
rect 108 748 180 836
rect 108 836 7236 924
<< m2 >>
rect 108 -44 7236 44
rect 7164 44 7236 132
rect 108 132 7092 220
rect 7164 132 7236 220
rect 108 220 180 308
rect 7164 220 7236 308
rect 108 308 180 396
rect 252 308 7236 396
rect 108 396 180 484
rect 7164 396 7236 484
rect 108 484 7092 572
rect 7164 484 7236 572
rect 108 572 180 660
rect 7164 572 7236 660
rect 108 660 180 748
rect 252 660 7236 748
rect 108 748 180 836
rect 108 836 7236 924
<< locali >>
rect 108 -44 7236 44
rect 7164 44 7236 132
rect 108 132 7092 220
rect 7164 132 7236 220
rect 108 220 180 308
rect 7164 220 7236 308
rect 108 308 180 396
rect 252 308 7236 396
rect 108 396 180 484
rect 7164 396 7236 484
rect 108 484 7092 572
rect 7164 484 7236 572
rect 108 572 180 660
rect 7164 572 7236 660
rect 108 660 180 748
rect 252 660 7236 748
rect 108 748 180 836
rect 108 836 7236 924
<< v1 >>
rect 6876 -35 6948 -26
rect 6876 -26 6948 -17
rect 6876 -17 6948 -8
rect 6876 -8 6948 0
rect 6876 0 6948 8
rect 6876 8 6948 17
rect 6876 17 6948 26
rect 6876 26 6948 35
rect 6948 -35 7020 -26
rect 6948 -26 7020 -17
rect 6948 -17 7020 -8
rect 6948 -8 7020 0
rect 6948 0 7020 8
rect 6948 8 7020 17
rect 6948 17 7020 26
rect 6948 26 7020 35
rect 7020 -35 7092 -26
rect 7020 -26 7092 -17
rect 7020 -17 7092 -8
rect 7020 -8 7092 0
rect 7020 0 7092 8
rect 7020 8 7092 17
rect 7020 17 7092 26
rect 7020 26 7092 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 6876 316 6948 325
rect 6876 325 6948 334
rect 6876 334 6948 343
rect 6876 343 6948 352
rect 6876 352 6948 360
rect 6876 360 6948 369
rect 6876 369 6948 378
rect 6876 378 6948 387
rect 6948 316 7020 325
rect 6948 325 7020 334
rect 6948 334 7020 343
rect 6948 343 7020 352
rect 6948 352 7020 360
rect 6948 360 7020 369
rect 6948 369 7020 378
rect 6948 378 7020 387
rect 7020 316 7092 325
rect 7020 325 7092 334
rect 7020 334 7092 343
rect 7020 343 7092 352
rect 7020 352 7092 360
rect 7020 360 7092 369
rect 7020 369 7092 378
rect 7020 378 7092 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 6876 668 6948 677
rect 6876 677 6948 686
rect 6876 686 6948 695
rect 6876 695 6948 704
rect 6876 704 6948 712
rect 6876 712 6948 721
rect 6876 721 6948 730
rect 6876 730 6948 739
rect 6948 668 7020 677
rect 6948 677 7020 686
rect 6948 686 7020 695
rect 6948 695 7020 704
rect 6948 704 7020 712
rect 6948 712 7020 721
rect 6948 721 7020 730
rect 6948 730 7020 739
rect 7020 668 7092 677
rect 7020 677 7092 686
rect 7020 686 7092 695
rect 7020 695 7092 704
rect 7020 704 7092 712
rect 7020 712 7092 721
rect 7020 721 7092 730
rect 7020 730 7092 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< v2 >>
rect 6876 -35 6948 -26
rect 6876 -26 6948 -17
rect 6876 -17 6948 -8
rect 6876 -8 6948 0
rect 6876 0 6948 8
rect 6876 8 6948 17
rect 6876 17 6948 26
rect 6876 26 6948 35
rect 6948 -35 7020 -26
rect 6948 -26 7020 -17
rect 6948 -17 7020 -8
rect 6948 -8 7020 0
rect 6948 0 7020 8
rect 6948 8 7020 17
rect 6948 17 7020 26
rect 6948 26 7020 35
rect 7020 -35 7092 -26
rect 7020 -26 7092 -17
rect 7020 -17 7092 -8
rect 7020 -8 7092 0
rect 7020 0 7092 8
rect 7020 8 7092 17
rect 7020 17 7092 26
rect 7020 26 7092 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 6876 316 6948 325
rect 6876 325 6948 334
rect 6876 334 6948 343
rect 6876 343 6948 352
rect 6876 352 6948 360
rect 6876 360 6948 369
rect 6876 369 6948 378
rect 6876 378 6948 387
rect 6948 316 7020 325
rect 6948 325 7020 334
rect 6948 334 7020 343
rect 6948 343 7020 352
rect 6948 352 7020 360
rect 6948 360 7020 369
rect 6948 369 7020 378
rect 6948 378 7020 387
rect 7020 316 7092 325
rect 7020 325 7092 334
rect 7020 334 7092 343
rect 7020 343 7092 352
rect 7020 352 7092 360
rect 7020 360 7092 369
rect 7020 369 7092 378
rect 7020 378 7092 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 6876 668 6948 677
rect 6876 677 6948 686
rect 6876 686 6948 695
rect 6876 695 6948 704
rect 6876 704 6948 712
rect 6876 712 6948 721
rect 6876 721 6948 730
rect 6876 730 6948 739
rect 6948 668 7020 677
rect 6948 677 7020 686
rect 6948 686 7020 695
rect 6948 695 7020 704
rect 6948 704 7020 712
rect 6948 712 7020 721
rect 6948 721 7020 730
rect 6948 730 7020 739
rect 7020 668 7092 677
rect 7020 677 7092 686
rect 7020 686 7092 695
rect 7020 695 7092 704
rect 7020 704 7092 712
rect 7020 712 7092 721
rect 7020 721 7092 730
rect 7020 730 7092 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< viali >>
rect 6876 -35 6948 -26
rect 6876 -26 6948 -17
rect 6876 -17 6948 -8
rect 6876 -8 6948 0
rect 6876 0 6948 8
rect 6876 8 6948 17
rect 6876 17 6948 26
rect 6876 26 6948 35
rect 6948 -35 7020 -26
rect 6948 -26 7020 -17
rect 6948 -17 7020 -8
rect 6948 -8 7020 0
rect 6948 0 7020 8
rect 6948 8 7020 17
rect 6948 17 7020 26
rect 6948 26 7020 35
rect 7020 -35 7092 -26
rect 7020 -26 7092 -17
rect 7020 -17 7092 -8
rect 7020 -8 7092 0
rect 7020 0 7092 8
rect 7020 8 7092 17
rect 7020 17 7092 26
rect 7020 26 7092 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 6876 316 6948 325
rect 6876 325 6948 334
rect 6876 334 6948 343
rect 6876 343 6948 352
rect 6876 352 6948 360
rect 6876 360 6948 369
rect 6876 369 6948 378
rect 6876 378 6948 387
rect 6948 316 7020 325
rect 6948 325 7020 334
rect 6948 334 7020 343
rect 6948 343 7020 352
rect 6948 352 7020 360
rect 6948 360 7020 369
rect 6948 369 7020 378
rect 6948 378 7020 387
rect 7020 316 7092 325
rect 7020 325 7092 334
rect 7020 334 7092 343
rect 7020 343 7092 352
rect 7020 352 7092 360
rect 7020 360 7092 369
rect 7020 369 7092 378
rect 7020 378 7092 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 6876 668 6948 677
rect 6876 677 6948 686
rect 6876 686 6948 695
rect 6876 695 6948 704
rect 6876 704 6948 712
rect 6876 712 6948 721
rect 6876 721 6948 730
rect 6876 730 6948 739
rect 6948 668 7020 677
rect 6948 677 7020 686
rect 6948 686 7020 695
rect 6948 695 7020 704
rect 6948 704 7020 712
rect 6948 712 7020 721
rect 6948 721 7020 730
rect 6948 730 7020 739
rect 7020 668 7092 677
rect 7020 677 7092 686
rect 7020 686 7092 695
rect 7020 695 7092 704
rect 7020 704 7092 712
rect 7020 712 7092 721
rect 7020 721 7092 730
rect 7020 730 7092 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< m3 >>
rect 108 -44 7236 44
rect 108 -44 7236 44
rect 7164 44 7236 132
rect 108 132 6876 220
rect 6948 132 7092 220
rect 7164 132 7236 220
rect 108 220 180 308
rect 7164 220 7236 308
rect 108 308 180 396
rect 252 308 324 396
rect 396 308 7236 396
rect 108 396 180 484
rect 7164 396 7236 484
rect 108 484 7092 572
rect 7164 484 7236 572
rect 108 572 180 660
rect 7164 572 7236 660
rect 108 660 180 748
rect 252 660 7236 748
rect 108 748 180 836
rect 108 836 7236 924
rect 108 836 7236 924
<< rm3 >>
rect 6876 132 6948 220
rect 324 308 396 396
<< labels >>
flabel m3 s 108 -44 7236 44 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 108 836 7236 924 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 7272 0 1056
<< end >>
