magic
tech sky130B
magscale 1 2
timestamp 1708642800
<< checkpaint >>
rect 0 0 2520 880
<< locali >>
rect 864 758 1032 826
rect 1032 54 1656 122
rect 1032 758 1656 826
rect 1032 54 1100 826
rect 398 142 466 738
rect 2054 142 2122 386
rect 2054 494 2122 738
rect 830 230 898 298
rect 830 406 898 474
rect 830 582 898 650
rect 1622 230 1690 298
rect 1622 406 1690 474
rect 1622 582 1690 650
rect 1980 142 2196 210
rect 1980 494 2196 562
rect 324 318 540 386
rect 756 758 972 826
rect 2412 132 2628 220
rect -108 132 108 220
<< m3 >>
rect 1548 0 1732 880
rect 756 0 940 880
rect 1548 0 1732 880
rect 756 0 940 880
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 176
box 0 176 1260 528
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_NCHDL MN3 
transform 1 0 0 0 1 528
box 0 528 1260 880
use SUNSAR_PCHDL MP0 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1 
transform 1 0 1260 0 1 176
box 1260 176 2520 528
use SUNSAR_PCHDL MP2 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_PCHDL MP3 
transform 1 0 1260 0 1 528
box 1260 528 2520 880
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 406
box 1548 406 1732 474
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 1548 0 1 406
box 1548 406 1732 474
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 756 0 1 54
box 756 54 940 122
use SUNSAR_cut_M1M4_2x1 xcut3 
transform 1 0 756 0 1 406
box 756 406 940 474
use SUNSAR_cut_M1M4_2x1 xcut4 
transform 1 0 756 0 1 406
box 756 406 940 474
<< labels >>
flabel locali s 1980 142 2196 210 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 1980 494 2196 562 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 324 318 540 386 0 FreeSans 400 0 0 0 RST
port 4 nsew signal bidirectional
flabel locali s 756 758 972 826 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 5 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 6 nsew signal bidirectional
flabel m3 s 1548 0 1732 880 0 FreeSans 400 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel m3 s 756 0 940 880 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 880
<< end >>
