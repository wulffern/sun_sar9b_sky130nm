magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect 0 0 7272 5280
<< m3 >>
rect -40 836 3672 912
rect -40 1892 3672 1968
rect -40 2948 3672 3024
rect -40 4004 3672 4080
rect -40 5060 3672 5136
rect -40 836 36 5136
rect 3672 -44 7308 32
rect 3672 1012 7308 1088
rect 3672 2068 7308 2144
rect 3672 3124 7308 3200
rect 3672 4180 7308 4256
rect 7308 -44 7384 4256
rect 108 2948 7236 3036
rect 108 -44 7236 44
use SUNSAR_CAP_BSSW_CV XCAPB0 
transform 1 0 0 0 1 0
box 0 0 7272 1056
use SUNSAR_CAP_BSSW_CV XCAPB1 
transform 1 0 0 0 1 1056
box 0 1056 7272 2112
use SUNSAR_CAP_BSSW_CV XCAPB2 
transform 1 0 0 0 1 2112
box 0 2112 7272 3168
use SUNSAR_CAP_BSSW_CV XCAPB3 
transform 1 0 0 0 1 3168
box 0 3168 7272 4224
use SUNSAR_CAP_BSSW_CV XCAPB4 
transform 1 0 0 0 1 4224
box 0 4224 7272 5280
<< labels >>
flabel m3 s 108 2948 7236 3036 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel m3 s 108 -44 7236 44 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 7272 0 5280
<< end >>
