magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 96 34
<< m3 >>
rect 0 0 92 34
<< v3 >>
rect 2 1 34 33
rect 58 1 90 33
<< m4 >>
rect 0 0 96 34
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 96 34
<< end >>
