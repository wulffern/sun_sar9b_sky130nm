magic
tech sky130B
magscale 1 2
timestamp 1708383600
<< checkpaint >>
rect 136 0 11404 27268
<< m1 >>
rect 2204 10332 2272 27200
rect 2204 10332 2272 27200
rect 2016 132 2084 27200
rect 2016 132 2084 27200
rect 1828 20532 1896 27200
rect 1828 20532 1896 27200
rect 1640 3532 1708 27200
rect 1640 3532 1708 27200
rect 1452 7536 1520 27200
rect 1452 7536 1520 27200
rect 1264 17736 1332 27200
rect 1264 17736 1332 27200
rect 1076 17132 1144 27200
rect 1076 17132 1144 27200
rect 888 18944 956 27200
rect 888 18944 956 27200
rect 700 8744 768 27200
rect 700 8744 768 27200
rect 512 9348 580 27200
rect 512 9348 580 27200
rect 324 8140 392 27200
rect 324 8140 392 27200
rect 136 9952 204 27200
rect 136 9952 204 27200
rect 2444 6932 2512 7116
rect 2444 6990 2756 7058
rect 2756 0 11336 68
<< m2 >>
rect 2272 10390 2444 10458
rect 2272 13410 2444 13478
rect 2272 11598 2444 11666
rect 2272 12806 2444 12874
rect 2272 12202 2444 12270
rect 2272 10994 2444 11062
rect 2272 23990 2444 24058
rect 2272 27010 2444 27078
rect 2272 25198 2444 25266
rect 2272 26406 2444 26474
rect 2272 25802 2444 25870
rect 2272 24594 2444 24662
rect 2084 190 2444 258
rect 2084 3210 2444 3278
rect 2084 1398 2444 1466
rect 2084 2606 2444 2674
rect 2084 2002 2444 2070
rect 2084 794 2444 862
rect 2084 13790 2444 13858
rect 2084 16810 2444 16878
rect 2084 14998 2444 15066
rect 2084 16206 2444 16274
rect 2084 15602 2444 15670
rect 2084 14394 2444 14462
rect 1896 20590 2444 20658
rect 1896 23610 2444 23678
rect 1896 21798 2444 21866
rect 1896 23006 2444 23074
rect 1896 22402 2444 22470
rect 1896 21194 2444 21262
rect 1708 3590 2444 3658
rect 1708 6610 2444 6678
rect 1708 4798 2444 4866
rect 1708 6006 2444 6074
rect 1708 5402 2444 5470
rect 1708 4194 2444 4262
rect 1520 7594 2444 7662
rect 1332 17794 2444 17862
rect 1144 17190 2444 17258
rect 1144 20210 2444 20278
rect 1144 18398 2444 18466
rect 1144 19606 2444 19674
rect 956 19002 2444 19070
rect 768 8802 2444 8870
rect 580 9406 2444 9474
rect 392 8198 2444 8266
rect 204 10010 2444 10078
<< locali >>
rect 2444 6932 2512 7116
<< viali >>
rect 2450 6944 2506 7000
rect 2450 7048 2506 7104
<< m3 >>
rect 2756 23800 2824 27268
use SUNSAR_CAP32C_CV XC1 
transform 1 0 2444 0 1 0
box 2444 0 11404 3400
use SUNSAR_CAP32C_CV XC64a<0> 
transform 1 0 2444 0 1 3400
box 2444 3400 11404 6800
use SUNSAR_CAP32C_CV XC32a<0> 
transform 1 0 2444 0 1 6800
box 2444 6800 11404 10200
use SUNSAR_CAP32C_CV XC128a<1> 
transform 1 0 2444 0 1 10200
box 2444 10200 11404 13600
use SUNSAR_CAP32C_CV XC128b<2> 
transform 1 0 2444 0 1 13600
box 2444 13600 11404 17000
use SUNSAR_CAP32C_CV X16ab 
transform 1 0 2444 0 1 17000
box 2444 17000 11404 20400
use SUNSAR_CAP32C_CV XC64b<1> 
transform 1 0 2444 0 1 20400
box 2444 20400 11404 23800
use SUNSAR_CAP32C_CV XC0 
transform 1 0 2444 0 1 23800
box 2444 23800 11404 27200
use SUNSAR_cut_M1M3_2x1 xcut0 
transform 1 0 2444 0 1 10390
box 2444 10390 2628 10458
use SUNSAR_cut_M2M3_1x2 xcut1 
transform 1 0 2204 0 1 10332
box 2204 10332 2272 10516
use SUNSAR_cut_M1M3_2x1 xcut2 
transform 1 0 2444 0 1 13410
box 2444 13410 2628 13478
use SUNSAR_cut_M2M3_1x2 xcut3 
transform 1 0 2204 0 1 13352
box 2204 13352 2272 13536
use SUNSAR_cut_M1M3_2x1 xcut4 
transform 1 0 2444 0 1 11598
box 2444 11598 2628 11666
use SUNSAR_cut_M2M3_1x2 xcut5 
transform 1 0 2204 0 1 11540
box 2204 11540 2272 11724
use SUNSAR_cut_M1M3_2x1 xcut6 
transform 1 0 2444 0 1 12806
box 2444 12806 2628 12874
use SUNSAR_cut_M2M3_1x2 xcut7 
transform 1 0 2204 0 1 12748
box 2204 12748 2272 12932
use SUNSAR_cut_M1M3_2x1 xcut8 
transform 1 0 2444 0 1 12202
box 2444 12202 2628 12270
use SUNSAR_cut_M2M3_1x2 xcut9 
transform 1 0 2204 0 1 12144
box 2204 12144 2272 12328
use SUNSAR_cut_M1M3_2x1 xcut10 
transform 1 0 2444 0 1 10994
box 2444 10994 2628 11062
use SUNSAR_cut_M2M3_1x2 xcut11 
transform 1 0 2204 0 1 10936
box 2204 10936 2272 11120
use SUNSAR_cut_M1M3_2x1 xcut12 
transform 1 0 2444 0 1 23990
box 2444 23990 2628 24058
use SUNSAR_cut_M2M3_1x2 xcut13 
transform 1 0 2204 0 1 23932
box 2204 23932 2272 24116
use SUNSAR_cut_M1M3_2x1 xcut14 
transform 1 0 2444 0 1 27010
box 2444 27010 2628 27078
use SUNSAR_cut_M2M3_1x2 xcut15 
transform 1 0 2204 0 1 26952
box 2204 26952 2272 27136
use SUNSAR_cut_M1M3_2x1 xcut16 
transform 1 0 2444 0 1 25198
box 2444 25198 2628 25266
use SUNSAR_cut_M2M3_1x2 xcut17 
transform 1 0 2204 0 1 25140
box 2204 25140 2272 25324
use SUNSAR_cut_M1M3_2x1 xcut18 
transform 1 0 2444 0 1 26406
box 2444 26406 2628 26474
use SUNSAR_cut_M2M3_1x2 xcut19 
transform 1 0 2204 0 1 26348
box 2204 26348 2272 26532
use SUNSAR_cut_M1M3_2x1 xcut20 
transform 1 0 2444 0 1 25802
box 2444 25802 2628 25870
use SUNSAR_cut_M2M3_1x2 xcut21 
transform 1 0 2204 0 1 25744
box 2204 25744 2272 25928
use SUNSAR_cut_M1M3_2x1 xcut22 
transform 1 0 2444 0 1 24594
box 2444 24594 2628 24662
use SUNSAR_cut_M2M3_1x2 xcut23 
transform 1 0 2204 0 1 24536
box 2204 24536 2272 24720
use SUNSAR_cut_M1M3_2x1 xcut24 
transform 1 0 2444 0 1 190
box 2444 190 2628 258
use SUNSAR_cut_M2M3_1x2 xcut25 
transform 1 0 2016 0 1 132
box 2016 132 2084 316
use SUNSAR_cut_M1M3_2x1 xcut26 
transform 1 0 2444 0 1 3210
box 2444 3210 2628 3278
use SUNSAR_cut_M2M3_1x2 xcut27 
transform 1 0 2016 0 1 3152
box 2016 3152 2084 3336
use SUNSAR_cut_M1M3_2x1 xcut28 
transform 1 0 2444 0 1 1398
box 2444 1398 2628 1466
use SUNSAR_cut_M2M3_1x2 xcut29 
transform 1 0 2016 0 1 1340
box 2016 1340 2084 1524
use SUNSAR_cut_M1M3_2x1 xcut30 
transform 1 0 2444 0 1 2606
box 2444 2606 2628 2674
use SUNSAR_cut_M2M3_1x2 xcut31 
transform 1 0 2016 0 1 2548
box 2016 2548 2084 2732
use SUNSAR_cut_M1M3_2x1 xcut32 
transform 1 0 2444 0 1 2002
box 2444 2002 2628 2070
use SUNSAR_cut_M2M3_1x2 xcut33 
transform 1 0 2016 0 1 1944
box 2016 1944 2084 2128
use SUNSAR_cut_M1M3_2x1 xcut34 
transform 1 0 2444 0 1 794
box 2444 794 2628 862
use SUNSAR_cut_M2M3_1x2 xcut35 
transform 1 0 2016 0 1 736
box 2016 736 2084 920
use SUNSAR_cut_M1M3_2x1 xcut36 
transform 1 0 2444 0 1 13790
box 2444 13790 2628 13858
use SUNSAR_cut_M2M3_1x2 xcut37 
transform 1 0 2016 0 1 13732
box 2016 13732 2084 13916
use SUNSAR_cut_M1M3_2x1 xcut38 
transform 1 0 2444 0 1 16810
box 2444 16810 2628 16878
use SUNSAR_cut_M2M3_1x2 xcut39 
transform 1 0 2016 0 1 16752
box 2016 16752 2084 16936
use SUNSAR_cut_M1M3_2x1 xcut40 
transform 1 0 2444 0 1 14998
box 2444 14998 2628 15066
use SUNSAR_cut_M2M3_1x2 xcut41 
transform 1 0 2016 0 1 14940
box 2016 14940 2084 15124
use SUNSAR_cut_M1M3_2x1 xcut42 
transform 1 0 2444 0 1 16206
box 2444 16206 2628 16274
use SUNSAR_cut_M2M3_1x2 xcut43 
transform 1 0 2016 0 1 16148
box 2016 16148 2084 16332
use SUNSAR_cut_M1M3_2x1 xcut44 
transform 1 0 2444 0 1 15602
box 2444 15602 2628 15670
use SUNSAR_cut_M2M3_1x2 xcut45 
transform 1 0 2016 0 1 15544
box 2016 15544 2084 15728
use SUNSAR_cut_M1M3_2x1 xcut46 
transform 1 0 2444 0 1 14394
box 2444 14394 2628 14462
use SUNSAR_cut_M2M3_1x2 xcut47 
transform 1 0 2016 0 1 14336
box 2016 14336 2084 14520
use SUNSAR_cut_M1M3_2x1 xcut48 
transform 1 0 2444 0 1 20590
box 2444 20590 2628 20658
use SUNSAR_cut_M2M3_1x2 xcut49 
transform 1 0 1828 0 1 20532
box 1828 20532 1896 20716
use SUNSAR_cut_M1M3_2x1 xcut50 
transform 1 0 2444 0 1 23610
box 2444 23610 2628 23678
use SUNSAR_cut_M2M3_1x2 xcut51 
transform 1 0 1828 0 1 23552
box 1828 23552 1896 23736
use SUNSAR_cut_M1M3_2x1 xcut52 
transform 1 0 2444 0 1 21798
box 2444 21798 2628 21866
use SUNSAR_cut_M2M3_1x2 xcut53 
transform 1 0 1828 0 1 21740
box 1828 21740 1896 21924
use SUNSAR_cut_M1M3_2x1 xcut54 
transform 1 0 2444 0 1 23006
box 2444 23006 2628 23074
use SUNSAR_cut_M2M3_1x2 xcut55 
transform 1 0 1828 0 1 22948
box 1828 22948 1896 23132
use SUNSAR_cut_M1M3_2x1 xcut56 
transform 1 0 2444 0 1 22402
box 2444 22402 2628 22470
use SUNSAR_cut_M2M3_1x2 xcut57 
transform 1 0 1828 0 1 22344
box 1828 22344 1896 22528
use SUNSAR_cut_M1M3_2x1 xcut58 
transform 1 0 2444 0 1 21194
box 2444 21194 2628 21262
use SUNSAR_cut_M2M3_1x2 xcut59 
transform 1 0 1828 0 1 21136
box 1828 21136 1896 21320
use SUNSAR_cut_M1M3_2x1 xcut60 
transform 1 0 2444 0 1 3590
box 2444 3590 2628 3658
use SUNSAR_cut_M2M3_1x2 xcut61 
transform 1 0 1640 0 1 3532
box 1640 3532 1708 3716
use SUNSAR_cut_M1M3_2x1 xcut62 
transform 1 0 2444 0 1 6610
box 2444 6610 2628 6678
use SUNSAR_cut_M2M3_1x2 xcut63 
transform 1 0 1640 0 1 6552
box 1640 6552 1708 6736
use SUNSAR_cut_M1M3_2x1 xcut64 
transform 1 0 2444 0 1 4798
box 2444 4798 2628 4866
use SUNSAR_cut_M2M3_1x2 xcut65 
transform 1 0 1640 0 1 4740
box 1640 4740 1708 4924
use SUNSAR_cut_M1M3_2x1 xcut66 
transform 1 0 2444 0 1 6006
box 2444 6006 2628 6074
use SUNSAR_cut_M2M3_1x2 xcut67 
transform 1 0 1640 0 1 5948
box 1640 5948 1708 6132
use SUNSAR_cut_M1M3_2x1 xcut68 
transform 1 0 2444 0 1 5402
box 2444 5402 2628 5470
use SUNSAR_cut_M2M3_1x2 xcut69 
transform 1 0 1640 0 1 5344
box 1640 5344 1708 5528
use SUNSAR_cut_M1M3_2x1 xcut70 
transform 1 0 2444 0 1 4194
box 2444 4194 2628 4262
use SUNSAR_cut_M2M3_1x2 xcut71 
transform 1 0 1640 0 1 4136
box 1640 4136 1708 4320
use SUNSAR_cut_M1M3_2x1 xcut72 
transform 1 0 2444 0 1 7594
box 2444 7594 2628 7662
use SUNSAR_cut_M2M3_1x2 xcut73 
transform 1 0 1452 0 1 7536
box 1452 7536 1520 7720
use SUNSAR_cut_M1M3_2x1 xcut74 
transform 1 0 2444 0 1 17794
box 2444 17794 2628 17862
use SUNSAR_cut_M2M3_1x2 xcut75 
transform 1 0 1264 0 1 17736
box 1264 17736 1332 17920
use SUNSAR_cut_M1M3_2x1 xcut76 
transform 1 0 2444 0 1 17190
box 2444 17190 2628 17258
use SUNSAR_cut_M2M3_1x2 xcut77 
transform 1 0 1076 0 1 17132
box 1076 17132 1144 17316
use SUNSAR_cut_M1M3_2x1 xcut78 
transform 1 0 2444 0 1 20210
box 2444 20210 2628 20278
use SUNSAR_cut_M2M3_1x2 xcut79 
transform 1 0 1076 0 1 20152
box 1076 20152 1144 20336
use SUNSAR_cut_M1M3_2x1 xcut80 
transform 1 0 2444 0 1 18398
box 2444 18398 2628 18466
use SUNSAR_cut_M2M3_1x2 xcut81 
transform 1 0 1076 0 1 18340
box 1076 18340 1144 18524
use SUNSAR_cut_M1M3_2x1 xcut82 
transform 1 0 2444 0 1 19606
box 2444 19606 2628 19674
use SUNSAR_cut_M2M3_1x2 xcut83 
transform 1 0 1076 0 1 19548
box 1076 19548 1144 19732
use SUNSAR_cut_M1M3_2x1 xcut84 
transform 1 0 2444 0 1 19002
box 2444 19002 2628 19070
use SUNSAR_cut_M2M3_1x2 xcut85 
transform 1 0 888 0 1 18944
box 888 18944 956 19128
use SUNSAR_cut_M1M3_2x1 xcut86 
transform 1 0 2444 0 1 8802
box 2444 8802 2628 8870
use SUNSAR_cut_M2M3_1x2 xcut87 
transform 1 0 700 0 1 8744
box 700 8744 768 8928
use SUNSAR_cut_M1M3_2x1 xcut88 
transform 1 0 2444 0 1 9406
box 2444 9406 2628 9474
use SUNSAR_cut_M2M3_1x2 xcut89 
transform 1 0 512 0 1 9348
box 512 9348 580 9532
use SUNSAR_cut_M1M3_2x1 xcut90 
transform 1 0 2444 0 1 8198
box 2444 8198 2628 8266
use SUNSAR_cut_M2M3_1x2 xcut91 
transform 1 0 324 0 1 8140
box 324 8140 392 8324
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 2444 0 1 10010
box 2444 10010 2628 10078
use SUNSAR_cut_M2M3_1x2 xcut93 
transform 1 0 136 0 1 9952
box 136 9952 204 10136
<< labels >>
flabel m1 s 2204 10332 2272 27200 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew signal bidirectional
flabel m1 s 2016 132 2084 27200 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew signal bidirectional
flabel m1 s 1828 20532 1896 27200 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew signal bidirectional
flabel m1 s 1640 3532 1708 27200 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew signal bidirectional
flabel m1 s 1452 7536 1520 27200 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew signal bidirectional
flabel m1 s 1264 17736 1332 27200 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew signal bidirectional
flabel m1 s 1076 17132 1144 27200 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew signal bidirectional
flabel m1 s 888 18944 956 27200 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew signal bidirectional
flabel m1 s 700 8744 768 27200 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew signal bidirectional
flabel m1 s 512 9348 580 27200 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew signal bidirectional
flabel m1 s 324 8140 392 27200 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew signal bidirectional
flabel m1 s 136 9952 204 27200 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew signal bidirectional
flabel m1 s 2756 0 11336 68 0 FreeSans 400 0 0 0 AVSS
port 14 nsew signal bidirectional
flabel m3 s 2756 23800 2824 27268 0 FreeSans 400 0 0 0 CTOP
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 136 11404 0 27268
<< end >>
