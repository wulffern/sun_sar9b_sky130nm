magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 34 92
<< m1 >>
rect 0 0 34 92
<< v1 >>
rect 3 6 31 34
rect 3 58 31 86
<< m2 >>
rect 0 0 34 92
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 34 92
<< end >>
