magic
tech sky130A
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 184 184
<< locali >>
rect 0 0 184 184
<< viali >>
rect 12 12 68 68
rect 12 116 68 172
rect 116 12 172 68
rect 116 116 172 172
<< m1 >>
rect 0 0 184 184
<< v1 >>
rect 12 12 68 68
rect 12 116 68 172
rect 116 12 172 68
rect 116 116 172 172
<< m2 >>
rect 0 0 184 184
<< v2 >>
rect 12 12 68 68
rect 12 116 68 172
rect 116 12 172 68
rect 116 116 172 172
<< m3 >>
rect 0 0 184 184
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 184 184
<< end >>
