magic
tech sky130A
timestamp 1713029161
<< poly >>
rect 162 79 1098 97
<< locali >>
rect 378 203 550 237
rect 162 159 270 193
rect 415 115 449 149
rect -54 66 54 110
rect 516 61 550 203
rect 912 159 1044 193
rect 774 115 882 149
rect 912 61 946 159
rect 990 71 1098 105
rect 1206 66 1314 110
rect 516 27 946 61
<< metal3 >>
rect 378 0 470 264
rect 774 0 866 264
use SUNSAR_NCHDL  MN0
timestamp 1712959200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_NCHDL  MN1
timestamp 1712959200
transform 1 0 0 0 1 88
box -90 -66 630 242
use SUNSAR_PCHDL  MP0
timestamp 1712959200
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_PCHDL  MP1
timestamp 1712959200
transform 1 0 630 0 1 88
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1712959200
transform 1 0 774 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1712959200
transform 1 0 378 0 1 27
box 0 0 92 34
<< labels >>
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 5 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 6 nsew signal bidirectional
flabel locali s 774 115 882 149 0 FreeSans 400 0 0 0 GNG
port 3 nsew signal bidirectional
flabel locali s 162 159 270 193 0 FreeSans 400 0 0 0 TIE_H
port 4 nsew signal bidirectional
flabel locali s 990 71 1098 105 0 FreeSans 400 0 0 0 C
port 1 nsew signal bidirectional
flabel locali s 378 203 486 237 0 FreeSans 400 0 0 0 GN
port 2 nsew signal bidirectional
flabel metal3 s 774 0 866 264 0 FreeSans 400 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel metal3 s 378 0 470 264 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 264
<< end >>
