magic
tech sky130A
timestamp 1712959200
<< checkpaint >>
rect 0 0 1260 440
<< poly >>
rect 162 343 1098 361
rect 162 255 1098 273
rect 162 167 1098 185
rect 162 79 1098 97
<< locali >>
rect -54 66 54 110
rect 199 105 233 369
rect 432 291 828 325
rect 516 149 550 291
rect 378 115 828 149
rect 162 71 270 105
rect 1027 71 1061 369
rect 1206 66 1314 110
<< metal3 >>
rect 378 0 470 440
rect 774 0 866 440
use SUNSAR_NCHDL  MN0
timestamp 1712959200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_NCHDL  MN1
timestamp 1712959200
transform 1 0 0 0 1 88
box -90 -66 630 242
use SUNSAR_NCHDL  MN2
timestamp 1712959200
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNSAR_NCHDL  MN3
timestamp 1712959200
transform 1 0 0 0 1 264
box -90 -66 630 242
use SUNSAR_PCHDL  MP0
timestamp 1712959200
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_PCHDL  MP1
timestamp 1712959200
transform 1 0 630 0 1 88
box 0 -66 720 242
use SUNSAR_PCHDL  MP2
timestamp 1712959200
transform 1 0 630 0 1 176
box 0 -66 720 242
use SUNSAR_PCHDL  MP3
timestamp 1712959200
transform 1 0 630 0 1 264
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1712959200
transform 1 0 774 0 1 27
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1712959200
transform 1 0 774 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut2
timestamp 1712959200
transform 1 0 774 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut3
timestamp 1712959200
transform 1 0 774 0 1 379
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut4
timestamp 1712959200
transform 1 0 378 0 1 27
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut5
timestamp 1712959200
transform 1 0 378 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut6
timestamp 1712959200
transform 1 0 378 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut7
timestamp 1712959200
transform 1 0 378 0 1 379
box 0 0 92 34
<< labels >>
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 378 115 486 149 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 3 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 4 nsew signal bidirectional
flabel metal3 s 774 0 866 440 0 FreeSans 400 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel metal3 s 378 0 470 440 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 440
<< end >>
