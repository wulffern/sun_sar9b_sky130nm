magic
tech sky130A
timestamp 1708968222
<< locali >>
rect 300 115 432 149
rect 828 115 946 149
rect 300 105 334 115
rect -54 71 334 105
rect 300 61 334 71
rect 912 105 946 115
rect 912 71 1314 105
rect 912 61 946 71
rect 300 27 432 61
rect 828 27 946 61
<< metal3 >>
rect 378 0 470 176
rect 774 0 866 176
use SUNSAR_NCHDL  MN1
timestamp 1708902000
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_PCHDL  MP1
timestamp 1708902000
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1708902000
transform 1 0 774 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1708902000
transform 1 0 774 0 1 27
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut2
timestamp 1708902000
transform 1 0 378 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut3
timestamp 1708902000
transform 1 0 378 0 1 27
box 0 0 92 34
<< labels >>
flabel metal3 s 774 0 866 176 0 FreeSans 200 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel metal3 s 378 0 470 176 0 FreeSans 200 0 0 0 AVSS
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
