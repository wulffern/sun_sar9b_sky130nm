magic
tech sky130B
magscale 1 2
timestamp 1672527600
<< checkpaint >>
rect 0 0 2520 1408
<< locali >>
rect 864 1290 1032 1350
rect 1032 58 1656 118
rect 1032 1290 1656 1350
rect 1032 58 1092 1350
rect 402 146 462 1262
rect 2058 146 2118 558
rect 2058 850 2118 1262
rect 834 234 894 470
rect 834 586 894 822
rect 834 938 894 1174
rect 1626 234 1686 470
rect 1626 586 1686 822
rect 1626 938 1686 1174
rect 1980 146 2196 206
rect 1980 850 2196 910
rect 324 498 540 558
rect 756 1290 972 1350
<< m3 >>
rect 1548 0 1748 1408
rect 756 0 956 1408
rect 1548 0 1748 1408
rect 756 0 956 1408
use SUNSAR_NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_NCHDL MN2
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNSAR_NCHDL MN3
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNSAR_PCHDL MP0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_PCHDL MP2
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNSAR_PCHDL MP3
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use SUNSAR_cut_M1M4_2x1 
transform 1 0 1548 0 1 586
box 1548 586 1748 662
use SUNSAR_cut_M1M4_2x1 
transform 1 0 1548 0 1 762
box 1548 762 1748 838
use SUNSAR_cut_M1M4_2x1 
transform 1 0 756 0 1 58
box 756 58 956 134
use SUNSAR_cut_M1M4_2x1 
transform 1 0 756 0 1 586
box 756 586 956 662
use SUNSAR_cut_M1M4_2x1 
transform 1 0 756 0 1 762
box 756 762 956 838
<< labels >>
flabel locali s 1980 146 2196 206 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 1980 850 2196 910 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 RST
port 4 nsew
flabel locali s 756 1290 972 1350 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel m3 s 1548 0 1748 1408 0 FreeSans 400 0 0 0 AVDD
port 7 nsew
flabel m3 s 756 0 956 1408 0 FreeSans 400 0 0 0 AVSS
port 8 nsew
<< end >>
