magic
tech sky130B
magscale 1 2
timestamp 1708642800
<< checkpaint >>
rect -1922 -1864 24278 37062
<< m3 >>
rect 8580 19144 22440 19212
rect 8580 19516 22440 19584
rect 20322 19856 20390 25540
rect 20598 19856 20666 30116
rect 194 19956 262 28708
rect 194 19956 262 28708
rect 4338 20142 4406 28708
rect 5234 20328 5302 28708
rect 884 20514 952 28738
rect 3763 20700 3831 28738
rect 3763 20700 3831 28738
rect 5924 20886 5992 28738
rect 5924 20886 5992 28738
rect 8803 21072 8871 28738
rect 8803 21072 8871 28738
rect 10964 21258 11032 28738
rect 10964 21258 11032 28738
rect 13843 21444 13911 28738
rect 13843 21444 13911 28738
rect 16004 21630 16072 28738
rect 16004 21630 16072 28738
rect 1027 21816 1095 29618
rect 3620 22002 3688 29618
rect 6067 22188 6135 29618
rect 1184 22374 1252 30498
rect 3464 22560 3532 30498
rect 6224 22746 6292 30498
rect 8504 22932 8572 30498
rect 11264 23118 11332 30498
rect 13544 23304 13612 30498
rect 16304 23490 16372 30498
rect 594 24166 778 35622
rect 3938 24166 4122 35622
rect 5634 24166 5818 35622
rect 8978 24166 9162 35622
rect 10674 24166 10858 35622
rect 14018 24166 14202 35622
rect 15714 24166 15898 35622
rect 19058 24166 19242 35622
rect 20754 24166 20938 35622
rect 8798 -720 8982 4800
rect 13374 -720 13558 4800
rect 1386 24166 1570 36342
rect 3146 24166 3330 36342
rect 6426 24166 6610 36342
rect 8186 24166 8370 36342
rect 11466 24166 11650 36342
rect 13226 24166 13410 36342
rect 16506 24166 16690 36342
rect 18266 24166 18450 36342
rect 21546 24166 21730 36342
rect 8006 -1440 8190 4800
rect 14166 -1440 14350 4800
rect 1962 28092 2146 37062
rect 2570 28092 2754 37062
rect 7002 28092 7186 37062
rect 7610 28092 7794 37062
rect 12042 28092 12226 37062
rect 12650 28092 12834 37062
rect 17082 28092 17266 37062
rect 17690 28092 17874 37062
rect 9376 -1864 9444 2938
rect 12912 -1864 12980 2938
rect 10078 1110 10314 1178
rect 8614 4986 10078 5054
rect 10078 1110 10146 5054
rect 12042 1110 12210 1178
rect 12210 4986 13742 5054
rect 12210 1110 12278 5054
rect 10314 1110 10482 1178
rect 10482 2518 12042 2586
rect 10482 1110 10550 2586
rect 10206 230 10390 298
rect 11966 230 12150 298
rect 18883 28738 18951 28922
<< m2 >>
rect 13708 18654 13776 19212
rect 8580 18654 8648 19584
rect 20322 19516 20390 19856
rect 20598 19144 20666 19856
rect 194 19888 13224 19956
rect 4338 20074 12848 20142
rect 5234 20260 12472 20328
rect 884 20446 9200 20514
rect 3763 20632 9576 20700
rect 5924 20818 9952 20886
rect 8803 21004 10328 21072
rect 10448 21190 11032 21258
rect 10636 21376 13911 21444
rect 10824 21562 16072 21630
rect 1027 21748 9388 21816
rect 3620 21934 9764 22002
rect 6067 22120 10140 22188
rect 1184 22306 13036 22374
rect 3464 22492 12660 22560
rect 6224 22678 12284 22746
rect 8504 22864 12096 22932
rect 11264 23050 11908 23118
rect 11652 23236 13612 23304
rect 11464 23422 16372 23490
rect 1386 34462 1722 34530
rect 1722 33860 4338 33928
rect 4270 33860 4338 34056
rect 1722 33860 1790 34530
rect 6426 34462 6762 34530
rect 6762 33860 9378 33928
rect 9310 33860 9378 34056
rect 6762 33860 6830 34530
rect 11466 34462 11802 34530
rect 11802 33860 14418 33928
rect 14350 33860 14418 34056
rect 11802 33860 11870 34530
rect 16506 34462 16842 34530
rect 16842 33860 19458 33928
rect 19390 33860 19458 34056
rect 16842 33860 16910 34530
rect 162 31396 19674 31464
rect 94 31396 162 31592
rect 4270 31396 4338 31592
rect 5134 31396 5202 31592
rect 9310 31396 9378 31592
rect 10174 31396 10242 31592
rect 14350 31396 14418 31592
rect 15214 31396 15282 31592
rect 19390 31396 19458 31592
rect 1418 24924 1722 24992
rect 1722 24532 4338 24600
rect 4270 24532 4338 24728
rect 1722 24532 1790 24992
rect 6458 24924 6762 24992
rect 6762 24532 9378 24600
rect 9310 24532 9378 24728
rect 6762 24532 6830 24992
rect 11498 24924 11802 24992
rect 11802 24532 14418 24600
rect 14350 24532 14418 24728
rect 11802 24532 11870 24992
rect 16538 24924 16842 24992
rect 16842 24532 19458 24600
rect 19390 24532 19458 24728
rect 16842 24532 16910 24992
rect 3114 24924 3418 24992
rect 3418 24924 3486 25052
rect 3418 25052 5234 25120
rect 5166 24660 5234 25120
rect 8154 24924 8458 24992
rect 8458 24924 8526 25052
rect 8458 25052 10274 25120
rect 10206 24660 10274 25120
rect 13194 24924 13498 24992
rect 13498 24924 13566 25052
rect 13498 25052 15314 25120
rect 15246 24660 15314 25120
rect 18234 24924 18538 24992
rect 18538 24924 18606 25052
rect 194 26696 19642 26764
rect 126 26420 194 26764
rect 4270 26420 4338 26764
rect 5166 26420 5234 26764
rect 9310 26420 9378 26764
rect 10206 26420 10274 26764
rect 14350 26420 14418 26764
rect 15246 26420 15314 26764
rect 19390 26420 19458 26764
rect 162 26848 19674 26916
rect 94 26848 162 27192
rect 4270 26848 4338 27192
rect 5134 26848 5202 27192
rect 9310 26848 9378 27192
rect 10174 26848 10242 27192
rect 14350 26848 14418 27192
rect 15214 26848 15282 27192
rect 19390 26848 19458 27192
rect 378 27476 1818 27544
rect 1818 27476 2898 27544
rect 1818 27476 7074 27544
rect 1818 27476 7938 27544
rect 1818 27476 12114 27544
rect 1818 27476 12978 27544
rect 1818 27476 17154 27544
rect 1818 27476 18018 27544
rect 702 32668 870 32736
rect 870 32668 938 32736
rect 4014 32668 4182 32736
rect 4182 32668 4250 32736
rect 5742 32668 5910 32736
rect 5910 32668 5978 32736
rect 9054 32668 9222 32736
rect 9222 32668 9290 32736
rect 10782 32668 10950 32736
rect 10950 32668 11018 32736
rect 14094 32668 14262 32736
rect 14262 32668 14330 32736
rect 15822 32668 15990 32736
rect 15990 32668 16058 32736
rect 19134 32668 19302 32736
rect 19302 33108 20430 33176
rect 19302 32668 19370 33176
rect 20206 27598 20862 27666
rect 19582 26488 20206 26556
rect 20206 26488 20274 27666
rect 19550 26420 19642 26488
rect 19566 27124 19734 27192
rect 19734 28512 21606 28580
rect 19734 27124 19802 28580
rect 21546 28444 21654 28512
rect 22086 32932 22254 33000
rect 19614 31808 22254 31876
rect 22254 31808 22322 33000
rect 19566 31876 19674 31944
rect 18342 34428 19866 34496
rect 19866 33494 20430 33562
rect 19866 33494 19934 34496
rect 10314 2518 10482 2586
rect 10482 1110 12042 1178
rect 10482 1110 10550 2586
rect 162 27476 2034 27544
<< m1 >>
rect 13156 18586 13224 19888
rect 12780 18586 12848 20074
rect 12404 18586 12472 20260
rect 9132 18586 9200 20446
rect 9508 18586 9576 20632
rect 9884 18586 9952 20818
rect 10260 18586 10328 21004
rect 10448 18586 10516 21190
rect 10636 18586 10704 21376
rect 10824 18586 10892 21562
rect 9320 18586 9388 21748
rect 9696 18586 9764 21934
rect 10072 18586 10140 22120
rect 12968 18586 13036 22306
rect 12592 18586 12660 22492
rect 12216 18586 12284 22678
rect 12028 18586 12096 22864
rect 11840 18586 11908 23050
rect 11652 18586 11720 23236
rect 11464 18586 11532 23422
rect 9272 -1652 9340 562
rect 13016 -1652 13084 562
rect -1854 33988 162 34056
rect 3114 34428 3450 34496
rect 3450 33860 5202 33928
rect 5134 33860 5202 34056
rect 3450 33860 3518 34496
rect 8154 34428 8490 34496
rect 8490 33860 10242 33928
rect 10174 33860 10242 34056
rect 8490 33860 8558 34496
rect 13194 34428 13530 34496
rect 13530 33860 15282 33928
rect 15214 33860 15282 34056
rect 13530 33860 13598 34496
rect -990 4986 68 5054
rect -990 8386 68 8454
rect -990 11786 68 11854
rect -990 15186 68 15254
rect 22288 4986 23346 5054
rect 22288 8386 23346 8454
rect 22288 11786 23346 11854
rect 22288 15186 23346 15254
<< locali >>
rect 23162 -720 23346 35622
rect -990 -720 23346 -536
rect -990 35438 23346 35622
rect -990 -720 -806 35622
rect 23162 -720 23346 35622
rect 23882 -1440 24066 36342
rect -1710 -1440 24066 -1256
rect -1710 36158 24066 36342
rect -1710 -1440 -1526 36342
rect 23882 -1440 24066 36342
rect -1710 36878 24066 37062
rect -1710 36878 24066 37062
rect 24210 -1652 24278 37062
rect -1710 -1652 24278 -1584
rect 24210 -1652 24278 37062
rect -1922 -1864 24278 -1796
rect -1922 -1864 -1854 37062
rect 19026 32668 19242 32736
rect 162 31524 378 31592
rect 1818 27476 2034 27544
rect 10206 2518 10422 2586
rect 10206 1110 10422 1178
use SUNSAR_SARBSSW_CV XB1 
transform -1 0 11178 0 1 0
box 11178 0 22626 4800
use SUNSAR_SARBSSW_CV XB2 
transform 1 0 11178 0 1 0
box 11178 0 22626 4800
use SUNSAR_CDAC7_CV XDAC1 
transform -1 0 11028 0 1 4986
box 11028 4986 21920 18654
use SUNSAR_CDAC7_CV XDAC2 
transform 1 0 11328 0 1 4986
box 11328 4986 22220 18654
use SUNSAR_SARDIGEX4_CV XA0 
transform 1 0 -162 0 1 24166
box -162 24166 2358 34902
use SUNSAR_SARDIGEX4_CV XA1 
transform -1 0 4878 0 1 24166
box 4878 24166 7398 34902
use SUNSAR_SARDIGEX4_CV XA2 
transform 1 0 4878 0 1 24166
box 4878 24166 7398 34902
use SUNSAR_SARDIGEX4_CV XA3 
transform -1 0 9918 0 1 24166
box 9918 24166 12438 34902
use SUNSAR_SARDIGEX4_CV XA4 
transform 1 0 9918 0 1 24166
box 9918 24166 12438 34902
use SUNSAR_SARDIGEX4_CV XA5 
transform -1 0 14958 0 1 24166
box 14958 24166 17478 34902
use SUNSAR_SARDIGEX4_CV XA6 
transform 1 0 14958 0 1 24166
box 14958 24166 17478 34902
use SUNSAR_SARDIGEX4_CV XA7 
transform -1 0 19998 0 1 24166
box 19998 24166 22518 34902
use SUNSAR_SARCMPX1_CV XA20 
transform 1 0 19998 0 1 24166
box 19998 24166 22518 34022
use SUNSAR_cut_M3M4_1x2 xcut0 
transform 1 0 13708 0 1 18654
box 13708 18654 13776 18838
use SUNSAR_cut_M3M4_2x1 xcut1 
transform 1 0 13708 0 1 19144
box 13708 19144 13892 19212
use SUNSAR_cut_M3M4_1x2 xcut2 
transform 1 0 8580 0 1 18654
box 8580 18654 8648 18838
use SUNSAR_cut_M3M4_2x1 xcut3 
transform 1 0 8580 0 1 19516
box 8580 19516 8764 19584
use SUNSAR_cut_M2M4_2x1 xcut4 
transform 1 0 20322 0 1 25540
box 20322 25540 20506 25608
use SUNSAR_cut_M3M4_2x1 xcut5 
transform 1 0 20322 0 1 19516
box 20322 19516 20506 19584
use SUNSAR_cut_M3M4_1x2 xcut6 
transform 1 0 20322 0 1 19856
box 20322 19856 20390 20040
use SUNSAR_cut_M3M4_2x1 xcut7 
transform 1 0 20482 0 1 30116
box 20482 30116 20666 30184
use SUNSAR_cut_M2M3_2x1 xcut8 
transform 1 0 20322 0 1 30116
box 20322 30116 20506 30184
use SUNSAR_cut_M3M4_2x1 xcut9 
transform 1 0 20598 0 1 19144
box 20598 19144 20782 19212
use SUNSAR_cut_M3M4_1x2 xcut10 
transform 1 0 20598 0 1 19856
box 20598 19856 20666 20040
use SUNSAR_cut_M3M4_1x2 xcut11 
transform 1 0 194 0 1 19830
box 194 19830 262 20014
use SUNSAR_cut_M2M3_1x2 xcut12 
transform 1 0 13156 0 1 19830
box 13156 19830 13224 20014
use SUNSAR_cut_M3M4_1x2 xcut13 
transform 1 0 4338 0 1 20016
box 4338 20016 4406 20200
use SUNSAR_cut_M2M3_1x2 xcut14 
transform 1 0 12780 0 1 20016
box 12780 20016 12848 20200
use SUNSAR_cut_M3M4_1x2 xcut15 
transform 1 0 5234 0 1 20202
box 5234 20202 5302 20386
use SUNSAR_cut_M2M3_1x2 xcut16 
transform 1 0 12404 0 1 20202
box 12404 20202 12472 20386
use SUNSAR_cut_M3M4_1x2 xcut17 
transform 1 0 884 0 1 20388
box 884 20388 952 20572
use SUNSAR_cut_M2M3_1x2 xcut18 
transform 1 0 9132 0 1 20388
box 9132 20388 9200 20572
use SUNSAR_cut_M3M4_1x2 xcut19 
transform 1 0 3763 0 1 20574
box 3763 20574 3831 20758
use SUNSAR_cut_M2M3_1x2 xcut20 
transform 1 0 9508 0 1 20574
box 9508 20574 9576 20758
use SUNSAR_cut_M3M4_1x2 xcut21 
transform 1 0 5924 0 1 20760
box 5924 20760 5992 20944
use SUNSAR_cut_M2M3_1x2 xcut22 
transform 1 0 9884 0 1 20760
box 9884 20760 9952 20944
use SUNSAR_cut_M3M4_1x2 xcut23 
transform 1 0 8803 0 1 20946
box 8803 20946 8871 21130
use SUNSAR_cut_M2M3_1x2 xcut24 
transform 1 0 10260 0 1 20946
box 10260 20946 10328 21130
use SUNSAR_cut_M3M4_1x2 xcut25 
transform 1 0 10964 0 1 21132
box 10964 21132 11032 21316
use SUNSAR_cut_M2M3_1x2 xcut26 
transform 1 0 10448 0 1 21132
box 10448 21132 10516 21316
use SUNSAR_cut_M3M4_1x2 xcut27 
transform 1 0 13843 0 1 21318
box 13843 21318 13911 21502
use SUNSAR_cut_M2M3_1x2 xcut28 
transform 1 0 10636 0 1 21318
box 10636 21318 10704 21502
use SUNSAR_cut_M3M4_1x2 xcut29 
transform 1 0 16004 0 1 21504
box 16004 21504 16072 21688
use SUNSAR_cut_M2M3_1x2 xcut30 
transform 1 0 10824 0 1 21504
box 10824 21504 10892 21688
use SUNSAR_cut_M3M4_1x2 xcut31 
transform 1 0 1027 0 1 21690
box 1027 21690 1095 21874
use SUNSAR_cut_M2M3_1x2 xcut32 
transform 1 0 9320 0 1 21690
box 9320 21690 9388 21874
use SUNSAR_cut_M3M4_1x2 xcut33 
transform 1 0 3620 0 1 21876
box 3620 21876 3688 22060
use SUNSAR_cut_M2M3_1x2 xcut34 
transform 1 0 9696 0 1 21876
box 9696 21876 9764 22060
use SUNSAR_cut_M3M4_1x2 xcut35 
transform 1 0 6067 0 1 22062
box 6067 22062 6135 22246
use SUNSAR_cut_M2M3_1x2 xcut36 
transform 1 0 10072 0 1 22062
box 10072 22062 10140 22246
use SUNSAR_cut_M3M4_1x2 xcut37 
transform 1 0 1184 0 1 22248
box 1184 22248 1252 22432
use SUNSAR_cut_M2M3_1x2 xcut38 
transform 1 0 12968 0 1 22248
box 12968 22248 13036 22432
use SUNSAR_cut_M3M4_1x2 xcut39 
transform 1 0 3464 0 1 22434
box 3464 22434 3532 22618
use SUNSAR_cut_M2M3_1x2 xcut40 
transform 1 0 12592 0 1 22434
box 12592 22434 12660 22618
use SUNSAR_cut_M3M4_1x2 xcut41 
transform 1 0 6224 0 1 22620
box 6224 22620 6292 22804
use SUNSAR_cut_M2M3_1x2 xcut42 
transform 1 0 12216 0 1 22620
box 12216 22620 12284 22804
use SUNSAR_cut_M3M4_1x2 xcut43 
transform 1 0 8504 0 1 22806
box 8504 22806 8572 22990
use SUNSAR_cut_M2M3_1x2 xcut44 
transform 1 0 12028 0 1 22806
box 12028 22806 12096 22990
use SUNSAR_cut_M3M4_1x2 xcut45 
transform 1 0 11264 0 1 22992
box 11264 22992 11332 23176
use SUNSAR_cut_M2M3_1x2 xcut46 
transform 1 0 11840 0 1 22992
box 11840 22992 11908 23176
use SUNSAR_cut_M3M4_1x2 xcut47 
transform 1 0 13544 0 1 23178
box 13544 23178 13612 23362
use SUNSAR_cut_M2M3_1x2 xcut48 
transform 1 0 11652 0 1 23178
box 11652 23178 11720 23362
use SUNSAR_cut_M3M4_1x2 xcut49 
transform 1 0 16304 0 1 23364
box 16304 23364 16372 23548
use SUNSAR_cut_M2M3_1x2 xcut50 
transform 1 0 11464 0 1 23364
box 11464 23364 11532 23548
use SUNSAR_cut_M1M4_2x2 xcut51 
transform 1 0 594 0 1 35438
box 594 35438 778 35622
use SUNSAR_cut_M1M4_2x2 xcut52 
transform 1 0 3938 0 1 35438
box 3938 35438 4122 35622
use SUNSAR_cut_M1M4_2x2 xcut53 
transform 1 0 5634 0 1 35438
box 5634 35438 5818 35622
use SUNSAR_cut_M1M4_2x2 xcut54 
transform 1 0 8978 0 1 35438
box 8978 35438 9162 35622
use SUNSAR_cut_M1M4_2x2 xcut55 
transform 1 0 10674 0 1 35438
box 10674 35438 10858 35622
use SUNSAR_cut_M1M4_2x2 xcut56 
transform 1 0 14018 0 1 35438
box 14018 35438 14202 35622
use SUNSAR_cut_M1M4_2x2 xcut57 
transform 1 0 15714 0 1 35438
box 15714 35438 15898 35622
use SUNSAR_cut_M1M4_2x2 xcut58 
transform 1 0 19058 0 1 35438
box 19058 35438 19242 35622
use SUNSAR_cut_M1M4_2x2 xcut59 
transform 1 0 20754 0 1 35438
box 20754 35438 20938 35622
use SUNSAR_cut_M1M4_2x2 xcut60 
transform 1 0 8798 0 1 -720
box 8798 -720 8982 -536
use SUNSAR_cut_M1M4_2x2 xcut61 
transform 1 0 13374 0 1 -720
box 13374 -720 13558 -536
use SUNSAR_cut_M1M4_2x2 xcut62 
transform 1 0 1386 0 1 36158
box 1386 36158 1570 36342
use SUNSAR_cut_M1M4_2x2 xcut63 
transform 1 0 3146 0 1 36158
box 3146 36158 3330 36342
use SUNSAR_cut_M1M4_2x2 xcut64 
transform 1 0 6426 0 1 36158
box 6426 36158 6610 36342
use SUNSAR_cut_M1M4_2x2 xcut65 
transform 1 0 8186 0 1 36158
box 8186 36158 8370 36342
use SUNSAR_cut_M1M4_2x2 xcut66 
transform 1 0 11466 0 1 36158
box 11466 36158 11650 36342
use SUNSAR_cut_M1M4_2x2 xcut67 
transform 1 0 13226 0 1 36158
box 13226 36158 13410 36342
use SUNSAR_cut_M1M4_2x2 xcut68 
transform 1 0 16506 0 1 36158
box 16506 36158 16690 36342
use SUNSAR_cut_M1M4_2x2 xcut69 
transform 1 0 18266 0 1 36158
box 18266 36158 18450 36342
use SUNSAR_cut_M1M4_2x2 xcut70 
transform 1 0 21546 0 1 36158
box 21546 36158 21730 36342
use SUNSAR_cut_M1M4_2x2 xcut71 
transform 1 0 8006 0 1 -1440
box 8006 -1440 8190 -1256
use SUNSAR_cut_M1M4_2x2 xcut72 
transform 1 0 14166 0 1 -1440
box 14166 -1440 14350 -1256
use SUNSAR_cut_M1M4_2x2 xcut73 
transform 1 0 1962 0 1 36878
box 1962 36878 2146 37062
use SUNSAR_cut_M1M4_2x2 xcut74 
transform 1 0 2570 0 1 36878
box 2570 36878 2754 37062
use SUNSAR_cut_M1M4_2x2 xcut75 
transform 1 0 7002 0 1 36878
box 7002 36878 7186 37062
use SUNSAR_cut_M1M4_2x2 xcut76 
transform 1 0 7610 0 1 36878
box 7610 36878 7794 37062
use SUNSAR_cut_M1M4_2x2 xcut77 
transform 1 0 12042 0 1 36878
box 12042 36878 12226 37062
use SUNSAR_cut_M1M4_2x2 xcut78 
transform 1 0 12650 0 1 36878
box 12650 36878 12834 37062
use SUNSAR_cut_M1M4_2x2 xcut79 
transform 1 0 17082 0 1 36878
box 17082 36878 17266 37062
use SUNSAR_cut_M1M4_2x2 xcut80 
transform 1 0 17690 0 1 36878
box 17690 36878 17874 37062
use SUNSAR_cut_M1M2_2x1 xcut81 
transform 1 0 9214 0 1 494
box 9214 494 9398 562
use SUNSAR_cut_M1M2_2x1 xcut82 
transform 1 0 9214 0 1 -1652
box 9214 -1652 9398 -1584
use SUNSAR_cut_M1M2_2x1 xcut83 
transform 1 0 12958 0 1 494
box 12958 494 13142 562
use SUNSAR_cut_M1M2_2x1 xcut84 
transform 1 0 12958 0 1 -1652
box 12958 -1652 13142 -1584
use SUNSAR_cut_M1M2_2x1 xcut85 
transform 1 0 162 0 1 33988
box 162 33988 346 34056
use SUNSAR_cut_M1M2_1x2 xcut86 
transform 1 0 -1922 0 1 33930
box -1922 33930 -1854 34114
use SUNSAR_cut_M1M4_2x1 xcut87 
transform 1 0 9318 0 1 -1864
box 9318 -1864 9502 -1796
use SUNSAR_cut_M1M4_2x1 xcut88 
transform 1 0 12854 0 1 -1864
box 12854 -1864 13038 -1796
use SUNSAR_cut_M1M3_2x1 xcut89 
transform 1 0 1386 0 1 34462
box 1386 34462 1570 34530
use SUNSAR_cut_M1M3_2x1 xcut90 
transform 1 0 4338 0 1 33988
box 4338 33988 4522 34056
use SUNSAR_cut_M1M3_2x1 xcut91 
transform 1 0 6426 0 1 34462
box 6426 34462 6610 34530
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 9378 0 1 33988
box 9378 33988 9562 34056
use SUNSAR_cut_M1M3_2x1 xcut93 
transform 1 0 11466 0 1 34462
box 11466 34462 11650 34530
use SUNSAR_cut_M1M3_2x1 xcut94 
transform 1 0 14418 0 1 33988
box 14418 33988 14602 34056
use SUNSAR_cut_M1M3_2x1 xcut95 
transform 1 0 16506 0 1 34462
box 16506 34462 16690 34530
use SUNSAR_cut_M1M3_2x1 xcut96 
transform 1 0 19458 0 1 33988
box 19458 33988 19642 34056
use SUNSAR_cut_M1M3_2x1 xcut97 
transform 1 0 162 0 1 31524
box 162 31524 346 31592
use SUNSAR_cut_M1M3_2x1 xcut98 
transform 1 0 4338 0 1 31524
box 4338 31524 4522 31592
use SUNSAR_cut_M1M3_2x1 xcut99 
transform 1 0 5202 0 1 31524
box 5202 31524 5386 31592
use SUNSAR_cut_M1M3_2x1 xcut100 
transform 1 0 9378 0 1 31524
box 9378 31524 9562 31592
use SUNSAR_cut_M1M3_2x1 xcut101 
transform 1 0 10242 0 1 31524
box 10242 31524 10426 31592
use SUNSAR_cut_M1M3_2x1 xcut102 
transform 1 0 14418 0 1 31524
box 14418 31524 14602 31592
use SUNSAR_cut_M1M3_2x1 xcut103 
transform 1 0 15282 0 1 31524
box 15282 31524 15466 31592
use SUNSAR_cut_M1M3_2x1 xcut104 
transform 1 0 19458 0 1 31524
box 19458 31524 19642 31592
use SUNSAR_cut_M1M2_2x1 xcut105 
transform 1 0 3114 0 1 34428
box 3114 34428 3298 34496
use SUNSAR_cut_M1M2_2x1 xcut106 
transform 1 0 5202 0 1 33988
box 5202 33988 5386 34056
use SUNSAR_cut_M1M2_2x1 xcut107 
transform 1 0 8154 0 1 34428
box 8154 34428 8338 34496
use SUNSAR_cut_M1M2_2x1 xcut108 
transform 1 0 10242 0 1 33988
box 10242 33988 10426 34056
use SUNSAR_cut_M1M2_2x1 xcut109 
transform 1 0 13194 0 1 34428
box 13194 34428 13378 34496
use SUNSAR_cut_M1M2_2x1 xcut110 
transform 1 0 15282 0 1 33988
box 15282 33988 15466 34056
use SUNSAR_cut_M1M3_2x1 xcut111 
transform 1 0 162 0 1 27124
box 162 27124 346 27192
use SUNSAR_cut_M1M3_2x1 xcut112 
transform 1 0 4338 0 1 27124
box 4338 27124 4522 27192
use SUNSAR_cut_M1M3_2x1 xcut113 
transform 1 0 5202 0 1 27124
box 5202 27124 5386 27192
use SUNSAR_cut_M1M3_2x1 xcut114 
transform 1 0 9378 0 1 27124
box 9378 27124 9562 27192
use SUNSAR_cut_M1M3_2x1 xcut115 
transform 1 0 10242 0 1 27124
box 10242 27124 10426 27192
use SUNSAR_cut_M1M3_2x1 xcut116 
transform 1 0 14418 0 1 27124
box 14418 27124 14602 27192
use SUNSAR_cut_M1M3_2x1 xcut117 
transform 1 0 15282 0 1 27124
box 15282 27124 15466 27192
use SUNSAR_cut_M1M3_2x1 xcut118 
transform 1 0 19458 0 1 27124
box 19458 27124 19642 27192
use SUNSAR_cut_M1M3_2x1 xcut119 
transform 1 0 1818 0 1 27476
box 1818 27476 2002 27544
use SUNSAR_cut_M1M3_2x1 xcut120 
transform 1 0 2682 0 1 27476
box 2682 27476 2866 27544
use SUNSAR_cut_M1M3_2x1 xcut121 
transform 1 0 6858 0 1 27476
box 6858 27476 7042 27544
use SUNSAR_cut_M1M3_2x1 xcut122 
transform 1 0 7722 0 1 27476
box 7722 27476 7906 27544
use SUNSAR_cut_M1M3_2x1 xcut123 
transform 1 0 11898 0 1 27476
box 11898 27476 12082 27544
use SUNSAR_cut_M1M3_2x1 xcut124 
transform 1 0 12762 0 1 27476
box 12762 27476 12946 27544
use SUNSAR_cut_M1M3_2x1 xcut125 
transform 1 0 16938 0 1 27476
box 16938 27476 17122 27544
use SUNSAR_cut_M1M3_2x1 xcut126 
transform 1 0 17802 0 1 27476
box 17802 27476 17986 27544
use SUNSAR_cut_M1M3_2x1 xcut127 
transform 1 0 594 0 1 32668
box 594 32668 778 32736
use SUNSAR_cut_M1M3_2x1 xcut128 
transform 1 0 3906 0 1 32668
box 3906 32668 4090 32736
use SUNSAR_cut_M1M3_2x1 xcut129 
transform 1 0 5634 0 1 32668
box 5634 32668 5818 32736
use SUNSAR_cut_M1M3_2x1 xcut130 
transform 1 0 8946 0 1 32668
box 8946 32668 9130 32736
use SUNSAR_cut_M1M3_2x1 xcut131 
transform 1 0 10674 0 1 32668
box 10674 32668 10858 32736
use SUNSAR_cut_M1M3_2x1 xcut132 
transform 1 0 13986 0 1 32668
box 13986 32668 14170 32736
use SUNSAR_cut_M1M3_2x1 xcut133 
transform 1 0 15714 0 1 32668
box 15714 32668 15898 32736
use SUNSAR_cut_M1M3_2x1 xcut134 
transform 1 0 19026 0 1 32668
box 19026 32668 19210 32736
use SUNSAR_cut_M1M3_2x1 xcut135 
transform 1 0 20322 0 1 33108
box 20322 33108 20506 33176
use SUNSAR_cut_M1M3_2x1 xcut136 
transform 1 0 20786 0 1 27598
box 20786 27598 20970 27666
use SUNSAR_cut_M1M3_2x1 xcut137 
transform 1 0 21546 0 1 28444
box 21546 28444 21730 28512
use SUNSAR_cut_M1M3_2x1 xcut138 
transform 1 0 21978 0 1 32932
box 21978 32932 22162 33000
use SUNSAR_cut_M1M3_2x1 xcut139 
transform 1 0 19458 0 1 31876
box 19458 31876 19642 31944
use SUNSAR_cut_M1M3_2x1 xcut140 
transform 1 0 18234 0 1 34428
box 18234 34428 18418 34496
use SUNSAR_cut_M1M3_2x1 xcut141 
transform 1 0 20322 0 1 33494
box 20322 33494 20506 33562
use SUNSAR_cut_M1M4_2x1 xcut142 
transform 1 0 11934 0 1 1110
box 11934 1110 12118 1178
use SUNSAR_cut_M1M3_2x1 xcut143 
transform 1 0 10206 0 1 2518
box 10206 2518 10390 2586
use SUNSAR_cut_M1M3_2x1 xcut144 
transform 1 0 11934 0 1 1110
box 11934 1110 12118 1178
use SUNSAR_cut_M1M4_2x1 xcut145 
transform 1 0 10206 0 1 1110
box 10206 1110 10390 1178
use SUNSAR_cut_M1M4_2x1 xcut146 
transform 1 0 11934 0 1 2518
box 11934 2518 12118 2586
use SUNSAR_cut_M1M3_2x1 xcut147 
transform 1 0 162 0 1 27476
box 162 27476 346 27544
use SUNSAR_cut_M1M2_2x2 xcut148 
transform 1 0 -990 0 1 5054
box -990 5054 -806 5238
use SUNSAR_cut_M1M2_2x2 xcut149 
transform 1 0 -990 0 1 8454
box -990 8454 -806 8638
use SUNSAR_cut_M1M2_2x2 xcut150 
transform 1 0 -990 0 1 11854
box -990 11854 -806 12038
use SUNSAR_cut_M1M2_2x2 xcut151 
transform 1 0 -990 0 1 15254
box -990 15254 -806 15438
use SUNSAR_cut_M1M2_1x2 xcut152 
transform 1 0 23278 0 1 4986
box 23278 4986 23346 5170
use SUNSAR_cut_M1M2_1x2 xcut153 
transform 1 0 23278 0 1 8386
box 23278 8386 23346 8570
use SUNSAR_cut_M1M2_1x2 xcut154 
transform 1 0 23278 0 1 11786
box 23278 11786 23346 11970
use SUNSAR_cut_M1M2_1x2 xcut155 
transform 1 0 23278 0 1 15186
box 23278 15186 23346 15370
<< labels >>
flabel m3 s 194 19956 262 28708 0 FreeSans 400 0 0 0 D<7>
port 6 nsew signal bidirectional
flabel m3 s 3763 20700 3831 28738 0 FreeSans 400 0 0 0 D<6>
port 7 nsew signal bidirectional
flabel m3 s 5924 20886 5992 28738 0 FreeSans 400 0 0 0 D<5>
port 8 nsew signal bidirectional
flabel m3 s 8803 21072 8871 28738 0 FreeSans 400 0 0 0 D<4>
port 9 nsew signal bidirectional
flabel m3 s 10964 21258 11032 28738 0 FreeSans 400 0 0 0 D<3>
port 10 nsew signal bidirectional
flabel m3 s 13843 21444 13911 28738 0 FreeSans 400 0 0 0 D<2>
port 11 nsew signal bidirectional
flabel m3 s 16004 21630 16072 28738 0 FreeSans 400 0 0 0 D<1>
port 12 nsew signal bidirectional
flabel locali s 23162 -720 23346 35622 0 FreeSans 400 0 0 0 AVSS
port 19 nsew signal bidirectional
flabel locali s 23882 -1440 24066 36342 0 FreeSans 400 0 0 0 AVDD
port 18 nsew signal bidirectional
flabel locali s -1710 36878 24066 37062 0 FreeSans 400 0 0 0 VREF
port 17 nsew signal bidirectional
flabel locali s 24210 -1652 24278 37062 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 16 nsew signal bidirectional
flabel locali s 19026 32668 19242 32736 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel m3 s 10206 230 10390 298 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel m3 s 11966 230 12150 298 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s 162 31524 378 31592 0 FreeSans 400 0 0 0 CK_SAMPLE
port 15 nsew signal bidirectional
flabel locali s 1818 27476 2034 27544 0 FreeSans 400 0 0 0 EN
port 14 nsew signal bidirectional
flabel locali s 10206 2518 10422 2586 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 10206 1110 10422 1178 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel m3 s 18883 28738 18951 28922 0 FreeSans 400 0 0 0 D<0>
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -1922 -1864 24278 37062
<< end >>
