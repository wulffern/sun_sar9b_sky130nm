magic
tech sky130B
magscale 1 2
timestamp 1680904800
<< checkpaint >>
rect 0 0 2520 1408
<< locali >>
rect 1626 586 1686 822
rect 1626 938 1686 1174
rect 864 234 1032 294
rect 864 586 1032 646
rect 864 762 1032 822
rect 1032 234 1092 822
rect 1428 410 1656 470
rect 864 1290 1428 1350
rect 1428 410 1488 1350
rect 1656 58 1824 118
rect 1824 1202 2088 1262
rect 1824 58 1884 1262
rect 756 58 1764 118
rect 2412 132 2628 220
rect -108 132 108 220
rect 324 850 540 910
rect 324 498 540 558
rect 1980 146 2196 206
rect 324 146 540 206
rect 1548 410 1764 470
<< poly >>
rect 324 510 2196 546
rect 324 862 2196 898
rect 324 1214 2196 1250
<< m3 >>
rect 1548 0 1748 1408
rect 756 0 956 1408
rect 1548 0 1748 1408
rect 756 0 956 1408
use SUNSAR_NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_NCHDL MN2
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNSAR_NCHDL MN3
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNSAR_PCHDL MP0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_PCHDL MP2
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNSAR_PCHDL MP3
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use SUNSAR_cut_M1M4_2x1 xcut0
transform 1 0 1548 0 1 234
box 1548 234 1748 310
use SUNSAR_cut_M1M4_2x1 xcut1
transform 1 0 1548 0 1 1290
box 1548 1290 1748 1366
use SUNSAR_cut_M1M4_2x1 xcut2
transform 1 0 756 0 1 410
box 756 410 956 486
use SUNSAR_cut_M1M4_2x1 xcut3
transform 1 0 756 0 1 938
box 756 938 956 1014
use SUNSAR_cut_M1M4_2x1 xcut4
transform 1 0 756 0 1 1114
box 756 1114 956 1190
<< labels >>
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel locali s 324 850 540 910 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 1980 146 2196 206 0 FreeSans 400 0 0 0 RST_N
port 5 nsew signal bidirectional
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 EN
port 3 nsew signal bidirectional
flabel locali s 1548 410 1764 470 0 FreeSans 400 0 0 0 ENO
port 4 nsew signal bidirectional
flabel m3 s 1548 0 1748 1408 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 756 0 956 1408 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 1408
<< end >>
