magic
tech sky130A
timestamp 1712959200
<< checkpaint >>
rect 0 0 1260 704
<< poly >>
rect 162 607 1098 625
rect 162 79 1098 97
<< locali >>
rect 378 643 744 677
rect 162 599 270 633
rect 710 589 744 643
rect 378 555 550 589
rect 199 193 233 545
rect 314 467 486 501
rect 314 325 348 467
rect 516 413 550 555
rect 415 379 550 413
rect 710 555 845 589
rect 710 413 744 555
rect 811 467 845 501
rect 1027 423 1061 633
rect 710 379 845 413
rect 314 291 449 325
rect 162 159 270 193
rect 314 149 348 291
rect 516 237 550 379
rect 1044 335 1162 369
rect 811 291 845 325
rect 415 203 845 237
rect 1128 193 1162 335
rect 1044 159 1162 193
rect 314 115 550 149
rect 811 115 845 149
rect -54 66 54 110
rect 162 71 270 105
rect 516 61 550 115
rect 1128 105 1162 159
rect 1044 71 1162 105
rect 1206 66 1314 110
rect 516 27 828 61
<< metal3 >>
rect 378 0 470 704
rect 774 325 866 704
rect 774 291 946 325
rect 774 0 866 291
rect 912 281 946 291
rect 912 247 1044 281
use SUNSAR_NCHDL  MN0
timestamp 1712959200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_NCHDL  MN1
timestamp 1712959200
transform 1 0 0 0 1 88
box -90 -66 630 242
use SUNSAR_NCHDL  MN2
timestamp 1712959200
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNSAR_NCHDL  MN3
timestamp 1712959200
transform 1 0 0 0 1 264
box -90 -66 630 242
use SUNSAR_NCHDL  MN4
timestamp 1712959200
transform 1 0 0 0 1 352
box -90 -66 630 242
use SUNSAR_NCHDL  MN5
timestamp 1712959200
transform 1 0 0 0 1 440
box -90 -66 630 242
use SUNSAR_NCHDL  MN6
timestamp 1712959200
transform 1 0 0 0 1 528
box -90 -66 630 242
use SUNSAR_PCHDL  MP0
timestamp 1712959200
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_PCHDL  MP1
timestamp 1712959200
transform 1 0 630 0 1 88
box 0 -66 720 242
use SUNSAR_PCHDL  MP2
timestamp 1712959200
transform 1 0 630 0 1 176
box 0 -66 720 242
use SUNSAR_PCHDL  MP3
timestamp 1712959200
transform 1 0 630 0 1 264
box 0 -66 720 242
use SUNSAR_PCHDL  MP4
timestamp 1712959200
transform 1 0 630 0 1 352
box 0 -66 720 242
use SUNSAR_PCHDL  MP5
timestamp 1712959200
transform 1 0 630 0 1 440
box 0 -66 720 242
use SUNSAR_PCHDL  MP6
timestamp 1712959200
transform 1 0 630 0 1 528
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1712959200
transform 1 0 774 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1712959200
transform 1 0 990 0 1 247
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut2
timestamp 1712959200
transform 1 0 774 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut3
timestamp 1712959200
transform 1 0 774 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut4
timestamp 1712959200
transform 1 0 774 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut5
timestamp 1712959200
transform 1 0 774 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut6
timestamp 1712959200
transform 1 0 774 0 1 467
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut7
timestamp 1712959200
transform 1 0 774 0 1 467
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut8
timestamp 1712959200
transform 1 0 774 0 1 643
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut9
timestamp 1712959200
transform 1 0 378 0 1 27
box 0 0 92 34
<< labels >>
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 7 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 8 nsew signal bidirectional
flabel locali s 378 467 486 501 0 FreeSans 400 0 0 0 N1
port 5 nsew signal bidirectional
flabel locali s 378 555 486 589 0 FreeSans 400 0 0 0 N2
port 6 nsew signal bidirectional
flabel locali s 162 159 270 193 0 FreeSans 400 0 0 0 CI
port 1 nsew signal bidirectional
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 378 643 486 677 0 FreeSans 400 0 0 0 CO
port 3 nsew signal bidirectional
flabel locali s 162 599 270 633 0 FreeSans 400 0 0 0 VMR
port 4 nsew signal bidirectional
flabel metal3 s 774 0 866 704 0 FreeSans 400 0 0 0 AVDD
port 9 nsew signal bidirectional
flabel metal3 s 378 0 470 704 0 FreeSans 400 0 0 0 AVSS
port 10 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 704
<< end >>
