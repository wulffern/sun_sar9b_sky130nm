magic
tech sky130A
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 2520 4224
<< locali >>
rect 1656 582 1824 650
rect 1824 954 2040 1022
rect 1824 582 1892 1022
rect 1980 1022 2088 1090
rect 1656 1110 1824 1178
rect 1824 1550 2088 1618
rect 1824 3662 2088 3730
rect 1824 1110 1892 3730
rect 432 2078 600 2146
rect 600 1110 864 1178
rect 600 1110 668 2146
rect 480 2890 600 2958
rect 600 1110 864 1178
rect 600 1110 668 2958
rect 432 2958 540 3026
rect 864 1638 1032 1706
rect 864 2166 1032 2234
rect 1032 1638 1100 2234
rect 432 4014 600 4082
rect 600 3750 864 3818
rect 600 3750 668 4082
rect 324 1374 540 1442
rect 324 494 540 562
rect 756 4102 972 4170
rect 756 3750 972 3818
rect 324 3310 540 3378
<< m1 >>
rect 2088 2078 2256 2146
rect 2088 2958 2256 3026
rect 1656 582 2256 650
rect 2256 582 2324 3026
rect 480 1482 600 1550
rect 600 758 864 826
rect 600 758 668 1550
rect 432 1550 540 1618
rect 480 3594 600 3662
rect 600 2890 2040 2958
rect 600 2890 668 3662
rect 432 3662 540 3730
rect 1980 2958 2088 3026
rect 864 3046 1032 3114
rect 864 3750 1032 3818
rect 1032 3046 1100 3818
rect 432 2430 600 2498
rect 600 2166 864 2234
rect 600 2166 668 2498
rect 1656 2518 1824 2586
rect 1824 1902 2088 1970
rect 1824 2782 2088 2850
rect 1824 1902 1892 2850
rect 1656 4102 1824 4170
rect 1824 3486 2088 3554
rect 1824 3486 1892 4170
rect 196 670 432 738
rect 196 3310 432 3378
rect 196 670 264 3378
<< m3 >>
rect 1548 0 1732 4224
rect 756 0 940 4224
rect 1548 0 1732 4224
rect 756 0 940 4224
use SUNSAR_TAPCELLB_CV XA0 
transform 1 0 0 0 1 0
box 0 0 2520 352
use SUNSAR_NDX1_CV XA1 
transform 1 0 0 0 1 352
box 0 352 2520 880
use SUNSAR_IVX1_CV XA2 
transform 1 0 0 0 1 880
box 0 880 2520 1232
use SUNSAR_IVTRIX1_CV XA3 
transform 1 0 0 0 1 1232
box 0 1232 2520 1760
use SUNSAR_IVTRIX1_CV XA4 
transform 1 0 0 0 1 1760
box 0 1760 2520 2288
use SUNSAR_IVX1_CV XA5 
transform 1 0 0 0 1 2288
box 0 2288 2520 2640
use SUNSAR_IVTRIX1_CV XA6 
transform 1 0 0 0 1 2640
box 0 2640 2520 3168
use SUNSAR_NDTRIX1_CV XA7 
transform 1 0 0 0 1 3168
box 0 3168 2520 3872
use SUNSAR_IVX1_CV XA8 
transform 1 0 0 0 1 3872
box 0 3872 2520 4224
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 1980 0 1 2078
box 1980 2078 2164 2146
use SUNSAR_cut_M1M2_2x1 xcut1 
transform 1 0 1980 0 1 2958
box 1980 2958 2164 3026
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 1548 0 1 582
box 1548 582 1732 650
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 324 0 1 1550
box 324 1550 508 1618
use SUNSAR_cut_M1M2_2x1 xcut4 
transform 1 0 756 0 1 758
box 756 758 940 826
use SUNSAR_cut_M1M2_2x1 xcut5 
transform 1 0 324 0 1 3662
box 324 3662 508 3730
use SUNSAR_cut_M1M2_2x1 xcut6 
transform 1 0 1980 0 1 2958
box 1980 2958 2164 3026
use SUNSAR_cut_M1M2_2x1 xcut7 
transform 1 0 756 0 1 3046
box 756 3046 940 3114
use SUNSAR_cut_M1M2_2x1 xcut8 
transform 1 0 756 0 1 3750
box 756 3750 940 3818
use SUNSAR_cut_M1M2_2x1 xcut9 
transform 1 0 324 0 1 2430
box 324 2430 508 2498
use SUNSAR_cut_M1M2_2x1 xcut10 
transform 1 0 756 0 1 2166
box 756 2166 940 2234
use SUNSAR_cut_M1M2_2x1 xcut11 
transform 1 0 1548 0 1 2518
box 1548 2518 1732 2586
use SUNSAR_cut_M1M2_2x1 xcut12 
transform 1 0 1980 0 1 1902
box 1980 1902 2164 1970
use SUNSAR_cut_M1M2_2x1 xcut13 
transform 1 0 1980 0 1 2782
box 1980 2782 2164 2850
use SUNSAR_cut_M1M2_2x1 xcut14 
transform 1 0 1548 0 1 4102
box 1548 4102 1732 4170
use SUNSAR_cut_M1M2_2x1 xcut15 
transform 1 0 1980 0 1 3486
box 1980 3486 2164 3554
use SUNSAR_cut_M1M2_2x1 xcut16 
transform 1 0 324 0 1 670
box 324 670 508 738
use SUNSAR_cut_M1M2_2x1 xcut17 
transform 1 0 324 0 1 3310
box 324 3310 508 3378
<< labels >>
flabel locali s 324 1374 540 1442 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 324 494 540 562 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 756 4102 972 4170 0 FreeSans 400 0 0 0 Q
port 4 nsew signal bidirectional
flabel locali s 756 3750 972 3818 0 FreeSans 400 0 0 0 QN
port 5 nsew signal bidirectional
flabel locali s 324 3310 540 3378 0 FreeSans 400 0 0 0 RN
port 3 nsew signal bidirectional
flabel m3 s 1548 0 1732 4224 0 FreeSans 400 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel m3 s 756 0 940 4224 0 FreeSans 400 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 4224
<< end >>
