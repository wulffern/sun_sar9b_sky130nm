magic
tech sky130A
timestamp 1712959200
<< checkpaint >>
rect 0 0 3636 480
<< locali >>
rect 54 416 3618 420
rect 54 384 162 416
rect 270 384 3618 416
rect 54 380 3618 384
rect 54 260 90 380
rect 126 336 3618 340
rect 126 304 3438 336
rect 3546 304 3618 336
rect 126 300 3618 304
rect 54 256 3546 260
rect 54 224 162 256
rect 270 224 3546 256
rect 54 220 3546 224
rect 54 100 90 220
rect 3582 180 3618 300
rect 126 176 3618 180
rect 126 144 3438 176
rect 3546 144 3618 176
rect 126 140 3618 144
rect 54 96 3546 100
rect 54 64 162 96
rect 270 64 3546 96
rect 54 60 3546 64
rect 3582 20 3618 140
rect 54 16 3618 20
rect 54 -16 3438 16
rect 3546 -16 3618 16
rect 54 -20 3618 -16
<< viali >>
rect 162 384 270 416
rect 3438 304 3546 336
rect 162 224 270 256
rect 3438 144 3546 176
rect 162 64 270 96
rect 3438 -16 3546 16
<< metal1 >>
rect 54 416 3618 420
rect 54 384 162 416
rect 270 384 3618 416
rect 54 380 3618 384
rect 54 260 90 380
rect 126 336 3618 340
rect 126 304 3438 336
rect 3546 304 3618 336
rect 126 300 3618 304
rect 54 256 3546 260
rect 54 224 162 256
rect 270 224 3546 256
rect 54 220 3546 224
rect 54 100 90 220
rect 3582 180 3618 300
rect 126 176 3618 180
rect 126 144 3438 176
rect 3546 144 3618 176
rect 126 140 3618 144
rect 54 96 3546 100
rect 54 64 162 96
rect 270 64 3546 96
rect 54 60 3546 64
rect 3582 20 3618 140
rect 54 16 3618 20
rect 54 -16 3438 16
rect 3546 -16 3618 16
rect 54 -20 3618 -16
<< via1 >>
rect 162 384 270 416
rect 3438 304 3546 336
rect 162 224 270 256
rect 3438 144 3546 176
rect 162 64 270 96
rect 3438 -16 3546 16
<< metal2 >>
rect 54 416 3618 420
rect 54 384 162 416
rect 270 384 3618 416
rect 54 380 3618 384
rect 54 260 90 380
rect 126 336 3618 340
rect 126 304 3438 336
rect 3546 304 3618 336
rect 126 300 3618 304
rect 54 256 3546 260
rect 54 224 162 256
rect 270 224 3546 256
rect 54 220 3546 224
rect 54 100 90 220
rect 3582 180 3618 300
rect 126 176 3618 180
rect 126 144 3438 176
rect 3546 144 3618 176
rect 126 140 3618 144
rect 54 96 3546 100
rect 54 64 162 96
rect 270 64 3546 96
rect 54 60 3546 64
rect 3582 20 3618 140
rect 54 16 3618 20
rect 54 -16 3438 16
rect 3546 -16 3618 16
rect 54 -20 3618 -16
<< via2 >>
rect 162 384 270 416
rect 3438 304 3546 336
rect 162 224 270 256
rect 3438 144 3546 176
rect 162 64 270 96
rect 3438 -16 3546 16
<< metal3 >>
rect 54 416 3618 420
rect 54 384 162 416
rect 270 384 3618 416
rect 54 380 3618 384
rect 54 260 90 380
rect 126 336 3618 340
rect 126 304 3438 336
rect 3546 304 3618 336
rect 126 300 3618 304
rect 54 256 3546 260
rect 54 224 162 256
rect 270 224 3546 256
rect 54 220 3546 224
rect 54 100 90 220
rect 3582 180 3618 300
rect 126 140 162 180
rect 198 176 3618 180
rect 198 144 3438 176
rect 3546 144 3618 176
rect 198 140 3618 144
rect 54 96 3438 100
rect 54 64 162 96
rect 270 64 3438 96
rect 54 60 3438 64
rect 3474 60 3546 100
rect 3582 20 3618 140
rect 54 16 3618 20
rect 54 -16 3438 16
rect 3546 -16 3618 16
rect 54 -20 3618 -16
<< rmetal3 >>
rect 162 140 198 180
rect 3438 60 3474 100
<< via3 >>
rect 162 384 270 416
rect 3438 304 3546 336
rect 162 224 270 256
rect 3438 144 3546 176
rect 162 64 270 96
rect 3438 -16 3546 16
<< metal4 >>
rect 54 416 3618 420
rect 54 384 162 416
rect 270 384 3618 416
rect 54 380 3618 384
rect 54 260 90 380
rect 126 336 3618 340
rect 126 304 3438 336
rect 3546 304 3618 336
rect 126 300 3618 304
rect 54 256 3546 260
rect 54 224 162 256
rect 270 224 3546 256
rect 54 220 3546 224
rect 54 100 90 220
rect 3582 180 3618 300
rect 126 176 3618 180
rect 126 144 3438 176
rect 3546 144 3618 176
rect 126 140 3618 144
rect 54 96 3546 100
rect 54 64 162 96
rect 270 64 3546 96
rect 54 60 3546 64
rect 3582 20 3618 140
rect 54 16 3618 20
rect 54 -16 3438 16
rect 3546 -16 3618 16
rect 54 -20 3618 -16
<< labels >>
flabel metal3 s 54 -20 3618 20 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel metal3 s 54 380 3618 420 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3636 480
<< end >>
