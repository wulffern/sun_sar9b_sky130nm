magic
tech sky130B
magscale 1 2
timestamp 1708642800
<< checkpaint >>
rect 0 0 2520 704
<< locali >>
rect 864 582 1032 650
rect 1032 582 1656 650
rect 1032 582 1100 650
rect 2054 142 2122 562
rect 830 230 898 298
rect 830 406 898 474
rect 1622 230 1690 298
rect 1622 406 1690 474
rect 2412 132 2628 220
rect -108 132 108 220
rect 324 142 540 210
rect 1980 494 2196 562
rect 324 494 540 562
rect 324 318 540 386
rect 756 582 972 650
<< m3 >>
rect 1548 0 1732 704
rect 756 0 940 704
rect 1548 0 1732 704
rect 756 0 940 704
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 176
box 0 176 1260 528
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_PCHDL MP0 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1 
transform 1 0 1260 0 1 176
box 1260 176 2520 528
use SUNSAR_PCHDL MP2 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 54
box 1548 54 1732 122
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 756 0 1 54
box 756 54 940 122
<< labels >>
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel locali s 324 142 540 210 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 1980 494 2196 562 0 FreeSans 400 0 0 0 RST_N
port 3 nsew signal bidirectional
flabel locali s 324 494 540 562 0 FreeSans 400 0 0 0 EN
port 4 nsew signal bidirectional
flabel locali s 324 318 540 386 0 FreeSans 400 0 0 0 LCK_N
port 5 nsew signal bidirectional
flabel locali s 756 582 972 650 0 FreeSans 400 0 0 0 CHL
port 2 nsew signal bidirectional
flabel m3 s 1548 0 1732 704 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 756 0 940 704 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 704
<< end >>
