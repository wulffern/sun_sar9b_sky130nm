magic
tech sky130B
magscale 1 2
timestamp 1708383600
<< checkpaint >>
rect 0 34 8960 3434
<< m3 >>
rect 312 0 380 3468
rect 312 0 380 3468
rect 444 132 512 3336
rect 576 0 644 3468
rect 708 132 776 3336
rect 840 0 908 3468
rect 972 132 1040 3336
rect 1104 0 1172 3468
rect 1236 132 1304 3336
rect 1368 0 1436 3468
rect 1500 132 1568 3336
rect 1632 0 1700 3468
rect 1764 132 1832 3336
rect 1896 0 1964 3468
rect 2028 132 2096 3336
rect 2160 0 2228 3468
rect 2292 132 2360 3336
rect 2424 0 2492 3468
rect 2556 132 2624 3336
rect 2688 0 2756 3468
rect 2820 132 2888 3336
rect 2952 0 3020 3468
rect 3084 132 3152 3336
rect 3216 0 3284 3468
rect 3348 132 3416 3336
rect 3480 0 3548 3468
rect 3612 132 3680 3336
rect 3744 0 3812 3468
rect 3876 132 3944 3336
rect 4008 0 4076 3468
rect 4140 132 4208 3336
rect 4272 0 4340 3468
rect 4404 132 4472 3336
rect 4536 0 4604 3468
rect 4668 132 4736 3336
rect 4800 0 4868 3468
rect 4932 132 5000 3336
rect 5064 0 5132 3468
rect 5196 132 5264 3336
rect 5328 0 5396 3468
rect 5460 132 5528 3336
rect 5592 0 5660 3468
rect 5724 132 5792 3336
rect 5856 0 5924 3468
rect 5988 132 6056 3336
rect 6120 0 6188 3468
rect 6252 132 6320 3336
rect 6384 0 6452 3468
rect 6516 132 6584 3336
rect 6648 0 6716 3468
rect 6780 132 6848 3336
rect 6912 0 6980 3468
rect 7044 132 7112 3336
rect 7176 0 7244 3468
rect 7308 132 7376 3336
rect 7440 0 7508 3468
rect 7572 132 7640 3336
rect 7704 0 7772 3468
rect 7836 132 7904 3336
rect 7968 0 8036 3468
rect 8100 132 8168 3336
rect 8232 0 8300 3468
rect 8364 132 8432 3336
rect 8496 0 8564 3468
rect 8628 132 8696 3336
rect 8892 0 8960 3468
rect 8760 0 8828 3468
rect 312 0 8760 68
rect 312 3400 8760 3468
<< m1 >>
rect 312 0 8892 68
rect 2292 376 2360 3468
rect 6780 0 6848 3092
rect 2556 0 2624 1280
rect 2556 1584 2624 3468
rect 6516 0 6584 1280
rect 6516 1584 6584 3468
rect 2028 0 2096 2488
rect 2028 2792 2096 3468
rect 2820 0 2888 2488
rect 2820 2792 2888 3468
rect 6252 0 6320 2488
rect 6252 2792 6320 3468
rect 7044 0 7112 2488
rect 7044 2792 7112 3468
rect 1500 0 1568 1884
rect 1500 2188 1568 3468
rect 1764 0 1832 1884
rect 1764 2188 1832 3468
rect 3084 0 3152 1884
rect 3084 2188 3152 3468
rect 3348 0 3416 1884
rect 3348 2188 3416 3468
rect 5724 0 5792 1884
rect 5724 2188 5792 3468
rect 5988 0 6056 1884
rect 5988 2188 6056 3468
rect 7308 0 7376 1884
rect 7308 2188 7376 3468
rect 7572 0 7640 1884
rect 7572 2188 7640 3468
rect 444 0 512 676
rect 444 980 512 3468
rect 708 0 776 676
rect 708 980 776 3468
rect 972 0 1040 676
rect 972 980 1040 3468
rect 1236 0 1304 676
rect 1236 980 1304 3468
rect 3612 0 3680 676
rect 3612 980 3680 3468
rect 3876 0 3944 676
rect 3876 980 3944 3468
rect 4140 0 4208 676
rect 4140 980 4208 3468
rect 4404 0 4472 676
rect 4404 980 4472 3468
rect 4668 0 4736 676
rect 4668 980 4736 3468
rect 4932 0 5000 676
rect 4932 980 5000 3468
rect 5196 0 5264 676
rect 5196 980 5264 3468
rect 5460 0 5528 676
rect 5460 980 5528 3468
rect 7836 0 7904 676
rect 7836 980 7904 3468
rect 8100 0 8168 676
rect 8100 980 8168 3468
rect 8364 0 8432 676
rect 8364 980 8432 3468
rect 8628 0 8696 676
rect 8628 980 8696 3468
rect 312 0 380 3400
rect 576 0 644 3400
rect 840 0 908 3400
rect 1104 0 1172 3400
rect 1368 0 1436 3400
rect 1632 0 1700 3400
rect 1896 0 1964 3400
rect 2160 0 2228 3400
rect 2424 0 2492 3400
rect 2688 0 2756 3400
rect 2952 0 3020 3400
rect 3216 0 3284 3400
rect 3480 0 3548 3400
rect 3744 0 3812 3400
rect 4008 0 4076 3400
rect 4272 0 4340 3400
rect 4536 0 4604 3400
rect 4800 0 4868 3400
rect 5064 0 5132 3400
rect 5328 0 5396 3400
rect 5592 0 5660 3400
rect 5856 0 5924 3400
rect 6120 0 6188 3400
rect 6384 0 6452 3400
rect 6648 0 6716 3400
rect 6912 0 6980 3400
rect 7176 0 7244 3400
rect 7440 0 7508 3400
rect 7704 0 7772 3400
rect 7968 0 8036 3400
rect 8232 0 8300 3400
rect 8496 0 8564 3400
rect 8892 0 8960 3468
rect 8760 0 8828 3468
rect 312 0 8892 68
rect 312 3400 8892 3468
<< locali >>
rect 0 190 184 258
rect 0 3210 184 3278
rect 0 1398 184 1466
rect 0 2606 184 2674
rect 0 2002 184 2070
rect 0 794 184 862
rect 320 794 8760 862
rect 320 190 8760 258
rect 320 3210 8760 3278
rect 320 1398 8760 1466
rect 320 2606 8760 2674
rect 320 2002 8760 2070
<< m2 >>
rect 8892 0 8960 3468
use SUNSAR_RM1 XRES1A 
transform 1 0 184 0 1 190
box 184 190 320 258
use SUNSAR_RM1 XRES1B 
transform 1 0 184 0 1 3210
box 184 3210 320 3278
use SUNSAR_RM1 XRES2 
transform 1 0 184 0 1 1398
box 184 1398 320 1466
use SUNSAR_RM1 XRES4 
transform 1 0 184 0 1 2606
box 184 2606 320 2674
use SUNSAR_RM1 XRES8 
transform 1 0 184 0 1 2002
box 184 2002 320 2070
use SUNSAR_RM1 XRES16 
transform 1 0 184 0 1 794
box 184 794 320 862
use SUNSAR_cut_M2M4_1x2 xcut0 
transform 1 0 8892 0 1 1550
box 8892 1550 8960 1734
use SUNSAR_cut_M1M4_1x2 xcut1 
transform 1 0 2292 0 1 132
box 2292 132 2360 316
use SUNSAR_cut_M1M4_1x2 xcut2 
transform 1 0 6780 0 1 3152
box 6780 3152 6848 3336
use SUNSAR_cut_M1M4_1x2 xcut3 
transform 1 0 2556 0 1 1340
box 2556 1340 2624 1524
use SUNSAR_cut_M1M4_1x2 xcut4 
transform 1 0 6516 0 1 1340
box 6516 1340 6584 1524
use SUNSAR_cut_M1M4_1x2 xcut5 
transform 1 0 2028 0 1 2548
box 2028 2548 2096 2732
use SUNSAR_cut_M1M4_1x2 xcut6 
transform 1 0 2820 0 1 2548
box 2820 2548 2888 2732
use SUNSAR_cut_M1M4_1x2 xcut7 
transform 1 0 6252 0 1 2548
box 6252 2548 6320 2732
use SUNSAR_cut_M1M4_1x2 xcut8 
transform 1 0 7044 0 1 2548
box 7044 2548 7112 2732
use SUNSAR_cut_M1M4_1x2 xcut9 
transform 1 0 1500 0 1 1944
box 1500 1944 1568 2128
use SUNSAR_cut_M1M4_1x2 xcut10 
transform 1 0 1764 0 1 1944
box 1764 1944 1832 2128
use SUNSAR_cut_M1M4_1x2 xcut11 
transform 1 0 3084 0 1 1944
box 3084 1944 3152 2128
use SUNSAR_cut_M1M4_1x2 xcut12 
transform 1 0 3348 0 1 1944
box 3348 1944 3416 2128
use SUNSAR_cut_M1M4_1x2 xcut13 
transform 1 0 5724 0 1 1944
box 5724 1944 5792 2128
use SUNSAR_cut_M1M4_1x2 xcut14 
transform 1 0 5988 0 1 1944
box 5988 1944 6056 2128
use SUNSAR_cut_M1M4_1x2 xcut15 
transform 1 0 7308 0 1 1944
box 7308 1944 7376 2128
use SUNSAR_cut_M1M4_1x2 xcut16 
transform 1 0 7572 0 1 1944
box 7572 1944 7640 2128
use SUNSAR_cut_M1M4_1x2 xcut17 
transform 1 0 444 0 1 736
box 444 736 512 920
use SUNSAR_cut_M1M4_1x2 xcut18 
transform 1 0 708 0 1 736
box 708 736 776 920
use SUNSAR_cut_M1M4_1x2 xcut19 
transform 1 0 972 0 1 736
box 972 736 1040 920
use SUNSAR_cut_M1M4_1x2 xcut20 
transform 1 0 1236 0 1 736
box 1236 736 1304 920
use SUNSAR_cut_M1M4_1x2 xcut21 
transform 1 0 3612 0 1 736
box 3612 736 3680 920
use SUNSAR_cut_M1M4_1x2 xcut22 
transform 1 0 3876 0 1 736
box 3876 736 3944 920
use SUNSAR_cut_M1M4_1x2 xcut23 
transform 1 0 4140 0 1 736
box 4140 736 4208 920
use SUNSAR_cut_M1M4_1x2 xcut24 
transform 1 0 4404 0 1 736
box 4404 736 4472 920
use SUNSAR_cut_M1M4_1x2 xcut25 
transform 1 0 4668 0 1 736
box 4668 736 4736 920
use SUNSAR_cut_M1M4_1x2 xcut26 
transform 1 0 4932 0 1 736
box 4932 736 5000 920
use SUNSAR_cut_M1M4_1x2 xcut27 
transform 1 0 5196 0 1 736
box 5196 736 5264 920
use SUNSAR_cut_M1M4_1x2 xcut28 
transform 1 0 5460 0 1 736
box 5460 736 5528 920
use SUNSAR_cut_M1M4_1x2 xcut29 
transform 1 0 7836 0 1 736
box 7836 736 7904 920
use SUNSAR_cut_M1M4_1x2 xcut30 
transform 1 0 8100 0 1 736
box 8100 736 8168 920
use SUNSAR_cut_M1M4_1x2 xcut31 
transform 1 0 8364 0 1 736
box 8364 736 8432 920
use SUNSAR_cut_M1M4_1x2 xcut32 
transform 1 0 8628 0 1 736
box 8628 736 8696 920
<< labels >>
flabel m3 s 312 0 380 3468 0 FreeSans 400 0 0 0 CTOP
port 7 nsew signal bidirectional
flabel m1 s 312 0 8892 68 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
flabel locali s 0 190 184 258 0 FreeSans 400 0 0 0 C1A
port 1 nsew signal bidirectional
flabel locali s 0 3210 184 3278 0 FreeSans 400 0 0 0 C1B
port 2 nsew signal bidirectional
flabel locali s 0 1398 184 1466 0 FreeSans 400 0 0 0 C2
port 3 nsew signal bidirectional
flabel locali s 0 2606 184 2674 0 FreeSans 400 0 0 0 C4
port 4 nsew signal bidirectional
flabel locali s 0 2002 184 2070 0 FreeSans 400 0 0 0 C8
port 5 nsew signal bidirectional
flabel locali s 0 794 184 862 0 FreeSans 400 0 0 0 C16
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 8960 34 3434
<< end >>
