magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect 0 0 200 76
<< m2 >>
rect 0 0 200 76
<< v2 >>
rect 12 6 76 70
rect 124 6 188 70
<< m3 >>
rect 0 0 200 76
<< labels >>
<< properties >>
string FIXED_BBOX 0 200 0 76
<< end >>
