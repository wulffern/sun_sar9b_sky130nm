magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect 0 0 11448 5280
<< m1 >>
rect 2988 1994 3420 2054
rect 3096 586 3264 646
rect 3264 850 3528 910
rect 3264 586 3324 910
rect 432 2610 600 2670
rect 600 3402 2304 3462
rect 600 2610 660 3462
rect 1872 2258 2040 2318
rect 2040 2728 3096 2788
rect 2040 2258 2100 2788
rect 864 938 1032 998
rect 1032 1642 2304 1702
rect 1032 938 1092 1702
<< locali >>
rect 636 234 864 294
rect 636 586 864 646
rect 636 938 864 998
rect 636 1290 864 1350
rect 636 1642 864 1702
rect 636 1994 864 2054
rect 636 2346 864 2406
rect 636 2698 864 2758
rect 636 234 696 2758
rect 402 146 462 1262
rect 402 1554 462 2670
rect 864 58 1032 118
rect 864 410 1032 470
rect 864 762 1032 822
rect 864 1114 1032 1174
rect 1032 58 1092 1174
rect 864 1466 1032 1526
rect 864 1818 1032 1878
rect 864 2170 1032 2230
rect 864 2522 1032 2582
rect 1032 1466 1092 2582
rect 1764 498 1980 558
rect 3420 850 3636 910
rect 756 1114 972 1174
rect 756 2522 972 2582
<< m2 >>
rect 1872 1906 2044 1982
rect 2044 616 2304 692
rect 2044 616 2120 1982
rect 1416 2346 2304 2422
rect 432 850 1416 926
rect 1416 850 1492 2422
rect 3096 1466 3268 1542
rect 3268 -44 4384 32
rect 3268 -44 3344 1542
<< m3 >>
rect 4136 2948 7848 3024
rect 3520 1994 4136 2070
rect 4136 1994 4212 3024
rect 772 226 972 302
rect 1612 3394 1812 3470
rect 2988 0 3188 5280
rect 2196 0 2396 5280
rect 2988 0 3188 5280
rect 2196 0 2396 5280
use SUNSAR_NCHDLR M1 
transform 1 0 0 0 1 0
box 0 0 1440 352
use SUNSAR_NCHDLR M2 
transform 1 0 0 0 1 352
box 0 352 1440 704
use SUNSAR_NCHDLR M3 
transform 1 0 0 0 1 704
box 0 704 1440 1056
use SUNSAR_NCHDLR M4 
transform 1 0 0 0 1 1056
box 0 1056 1440 1408
use SUNSAR_NCHDLR M5 
transform 1 0 0 0 1 1408
box 0 1408 1440 1760
use SUNSAR_NCHDLR M6 
transform 1 0 0 0 1 1760
box 0 1760 1440 2112
use SUNSAR_NCHDLR M7 
transform 1 0 0 0 1 2112
box 0 2112 1440 2464
use SUNSAR_NCHDLR M8 
transform 1 0 0 0 1 2464
box 0 2464 1440 2816
use SUNSAR_TAPCELLB_CV XA5b 
transform 1 0 1440 0 1 0
box 1440 0 3960 352
use SUNSAR_IVX1_CV XA0 
transform 1 0 1440 0 1 352
box 1440 352 3960 704
use SUNSAR_TGPD_CV XA3 
transform 1 0 1440 0 1 704
box 1440 704 3960 1760
use SUNSAR_SARBSSWCTRL_CV XA4 
transform 1 0 1440 0 1 1760
box 1440 1760 3960 2464
use SUNSAR_TIEH_CV XA1 
transform 1 0 1440 0 1 2464
box 1440 2464 3960 2816
use SUNSAR_TAPCELLB_CV XA7 
transform 1 0 1440 0 1 2816
box 1440 2816 3960 3168
use SUNSAR_TIEL_CV XA2 
transform 1 0 1440 0 1 3168
box 1440 3168 3960 3520
use SUNSAR_TAPCELLB_CV XA5 
transform 1 0 1440 0 1 3520
box 1440 3520 3960 3872
use SUNSAR_CAP_BSSW5_CV XCAPB1 
transform 1 0 4176 0 1 0
box 4176 0 11448 5280
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 2988 0 1 1994
box 2988 1994 3172 2062
use SUNSAR_cut_M2M4_2x1 xcut1 
transform 1 0 3420 0 1 1994
box 3420 1994 3620 2070
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 2988 0 1 586
box 2988 586 3172 654
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 3420 0 1 850
box 3420 850 3604 918
use SUNSAR_cut_M1M3_2x1 xcut4 
transform 1 0 1764 0 1 1906
box 1764 1906 1964 1982
use SUNSAR_cut_M1M3_2x1 xcut5 
transform 1 0 2196 0 1 624
box 2196 624 2396 700
use SUNSAR_cut_M1M2_2x1 xcut6 
transform 1 0 324 0 1 2610
box 324 2610 508 2678
use SUNSAR_cut_M1M2_2x1 xcut7 
transform 1 0 2196 0 1 3402
box 2196 3402 2380 3470
use SUNSAR_cut_M1M2_2x1 xcut8 
transform 1 0 1764 0 1 2258
box 1764 2258 1948 2326
use SUNSAR_cut_M1M2_2x1 xcut9 
transform 1 0 2988 0 1 2732
box 2988 2732 3172 2800
use SUNSAR_cut_M1M2_2x1 xcut10 
transform 1 0 756 0 1 938
box 756 938 940 1006
use SUNSAR_cut_M1M2_2x1 xcut11 
transform 1 0 2196 0 1 1642
box 2196 1642 2380 1710
use SUNSAR_cut_M1M3_2x1 xcut12 
transform 1 0 2212 0 1 2346
box 2212 2346 2412 2422
use SUNSAR_cut_M1M3_2x1 xcut13 
transform 1 0 340 0 1 850
box 340 850 540 926
use SUNSAR_cut_M1M3_2x1 xcut14 
transform 1 0 2988 0 1 1466
box 2988 1466 3188 1542
use SUNSAR_cut_M3M4_2x1 xcut15 
transform 1 0 4284 0 1 -44
box 4284 -44 4484 32
use SUNSAR_cut_M1M4_2x1 xcut16 
transform 1 0 772 0 1 226
box 772 226 972 302
use SUNSAR_cut_M2M4_2x1 xcut17 
transform 1 0 1612 0 1 3394
box 1612 3394 1812 3470
<< labels >>
flabel m3 s 772 226 972 302 0 FreeSans 400 0 0 0 VI
port 1 nsew signal bidirectional
flabel m3 s 1612 3394 1812 3470 0 FreeSans 400 0 0 0 TIE_L
port 4 nsew signal bidirectional
flabel locali s 1764 498 1980 558 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 3420 850 3636 910 0 FreeSans 400 0 0 0 CKN
port 3 nsew signal bidirectional
flabel locali s 756 1114 972 1174 0 FreeSans 400 0 0 0 VO1
port 5 nsew signal bidirectional
flabel locali s 756 2522 972 2582 0 FreeSans 400 0 0 0 VO2
port 6 nsew signal bidirectional
flabel m3 s 2988 0 3188 5280 0 FreeSans 400 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel m3 s 2196 0 2396 5280 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 11448 0 5280
<< end >>
