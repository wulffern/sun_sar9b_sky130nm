magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 68 0 5974 13922
<< m1 >>
rect 1102 5282 1136 13888
rect 1102 5282 1136 13888
rect 1008 74 1042 13888
rect 1008 74 1042 13888
rect 914 10490 948 13888
rect 914 10490 948 13888
rect 820 1810 854 13888
rect 820 1810 854 13888
rect 726 3852 760 13888
rect 726 3852 760 13888
rect 632 9060 666 13888
rect 632 9060 666 13888
rect 538 8754 572 13888
rect 538 8754 572 13888
rect 444 9672 478 13888
rect 444 9672 478 13888
rect 350 4464 384 13888
rect 350 4464 384 13888
rect 256 4770 290 13888
rect 256 4770 290 13888
rect 162 4158 196 13888
rect 162 4158 196 13888
rect 68 5076 102 13888
rect 68 5076 102 13888
rect 1222 3546 1256 3638
rect 1222 3573 1386 3607
rect 1386 0 5936 38
<< m2 >>
rect 1136 5309 1222 5347
rect 1136 6839 1222 6877
rect 1136 5921 1222 5959
rect 1136 6533 1222 6571
rect 1136 6227 1222 6265
rect 1136 5615 1222 5653
rect 1136 12253 1222 12291
rect 1136 13783 1222 13821
rect 1136 12865 1222 12903
rect 1136 13477 1222 13515
rect 1136 13171 1222 13209
rect 1136 12559 1222 12597
rect 1042 101 1222 139
rect 1042 1631 1222 1669
rect 1042 713 1222 751
rect 1042 1325 1222 1363
rect 1042 1019 1222 1057
rect 1042 407 1222 445
rect 1042 7045 1222 7083
rect 1042 8575 1222 8613
rect 1042 7657 1222 7695
rect 1042 8269 1222 8307
rect 1042 7963 1222 8001
rect 1042 7351 1222 7389
rect 948 10517 1222 10555
rect 948 12047 1222 12085
rect 948 11129 1222 11167
rect 948 11741 1222 11779
rect 948 11435 1222 11473
rect 948 10823 1222 10861
rect 854 1837 1222 1875
rect 854 3367 1222 3405
rect 854 2449 1222 2487
rect 854 3061 1222 3099
rect 854 2755 1222 2793
rect 854 2143 1222 2181
rect 760 3879 1222 3917
rect 666 9087 1222 9125
rect 572 8781 1222 8819
rect 572 10311 1222 10349
rect 572 9393 1222 9431
rect 572 10005 1222 10043
rect 478 9699 1222 9737
rect 384 4491 1222 4529
rect 290 4797 1222 4835
rect 196 4185 1222 4223
rect 102 5103 1222 5141
<< locali >>
rect 1222 3546 1256 3638
<< viali >>
rect 1225 3552 1253 3580
rect 1225 3604 1253 3632
<< m3 >>
rect 1386 12152 1424 13922
use SUNSAR_CAP32C_CV XC1 
transform 1 0 1222 0 1 0
box 1222 0 5974 1736
use SUNSAR_CAP32C_CV XC64a<0> 
transform 1 0 1222 0 1 1736
box 1222 1736 5974 3472
use SUNSAR_CAP32C_CV XC32a<0> 
transform 1 0 1222 0 1 3472
box 1222 3472 5974 5208
use SUNSAR_CAP32C_CV XC128a<1> 
transform 1 0 1222 0 1 5208
box 1222 5208 5974 6944
use SUNSAR_CAP32C_CV XC128b<2> 
transform 1 0 1222 0 1 6944
box 1222 6944 5974 8680
use SUNSAR_CAP32C_CV X16ab 
transform 1 0 1222 0 1 8680
box 1222 8680 5974 10416
use SUNSAR_CAP32C_CV XC64b<1> 
transform 1 0 1222 0 1 10416
box 1222 10416 5974 12152
use SUNSAR_CAP32C_CV XC0 
transform 1 0 1222 0 1 12152
box 1222 12152 5974 13888
use SUNSAR_cut_M1M3_2x1 xcut0 
transform 1 0 1222 0 1 5309
box 1222 5309 1314 5343
use SUNSAR_cut_M2M3_1x2 xcut1 
transform 1 0 1102 0 1 5282
box 1102 5282 1136 5374
use SUNSAR_cut_M1M3_2x1 xcut2 
transform 1 0 1222 0 1 6839
box 1222 6839 1314 6873
use SUNSAR_cut_M2M3_1x2 xcut3 
transform 1 0 1102 0 1 6812
box 1102 6812 1136 6904
use SUNSAR_cut_M1M3_2x1 xcut4 
transform 1 0 1222 0 1 5921
box 1222 5921 1314 5955
use SUNSAR_cut_M2M3_1x2 xcut5 
transform 1 0 1102 0 1 5894
box 1102 5894 1136 5986
use SUNSAR_cut_M1M3_2x1 xcut6 
transform 1 0 1222 0 1 6533
box 1222 6533 1314 6567
use SUNSAR_cut_M2M3_1x2 xcut7 
transform 1 0 1102 0 1 6506
box 1102 6506 1136 6598
use SUNSAR_cut_M1M3_2x1 xcut8 
transform 1 0 1222 0 1 6227
box 1222 6227 1314 6261
use SUNSAR_cut_M2M3_1x2 xcut9 
transform 1 0 1102 0 1 6200
box 1102 6200 1136 6292
use SUNSAR_cut_M1M3_2x1 xcut10 
transform 1 0 1222 0 1 5615
box 1222 5615 1314 5649
use SUNSAR_cut_M2M3_1x2 xcut11 
transform 1 0 1102 0 1 5588
box 1102 5588 1136 5680
use SUNSAR_cut_M1M3_2x1 xcut12 
transform 1 0 1222 0 1 12253
box 1222 12253 1314 12287
use SUNSAR_cut_M2M3_1x2 xcut13 
transform 1 0 1102 0 1 12226
box 1102 12226 1136 12318
use SUNSAR_cut_M1M3_2x1 xcut14 
transform 1 0 1222 0 1 13783
box 1222 13783 1314 13817
use SUNSAR_cut_M2M3_1x2 xcut15 
transform 1 0 1102 0 1 13756
box 1102 13756 1136 13848
use SUNSAR_cut_M1M3_2x1 xcut16 
transform 1 0 1222 0 1 12865
box 1222 12865 1314 12899
use SUNSAR_cut_M2M3_1x2 xcut17 
transform 1 0 1102 0 1 12838
box 1102 12838 1136 12930
use SUNSAR_cut_M1M3_2x1 xcut18 
transform 1 0 1222 0 1 13477
box 1222 13477 1314 13511
use SUNSAR_cut_M2M3_1x2 xcut19 
transform 1 0 1102 0 1 13450
box 1102 13450 1136 13542
use SUNSAR_cut_M1M3_2x1 xcut20 
transform 1 0 1222 0 1 13171
box 1222 13171 1314 13205
use SUNSAR_cut_M2M3_1x2 xcut21 
transform 1 0 1102 0 1 13144
box 1102 13144 1136 13236
use SUNSAR_cut_M1M3_2x1 xcut22 
transform 1 0 1222 0 1 12559
box 1222 12559 1314 12593
use SUNSAR_cut_M2M3_1x2 xcut23 
transform 1 0 1102 0 1 12532
box 1102 12532 1136 12624
use SUNSAR_cut_M1M3_2x1 xcut24 
transform 1 0 1222 0 1 101
box 1222 101 1314 135
use SUNSAR_cut_M2M3_1x2 xcut25 
transform 1 0 1008 0 1 74
box 1008 74 1042 166
use SUNSAR_cut_M1M3_2x1 xcut26 
transform 1 0 1222 0 1 1631
box 1222 1631 1314 1665
use SUNSAR_cut_M2M3_1x2 xcut27 
transform 1 0 1008 0 1 1604
box 1008 1604 1042 1696
use SUNSAR_cut_M1M3_2x1 xcut28 
transform 1 0 1222 0 1 713
box 1222 713 1314 747
use SUNSAR_cut_M2M3_1x2 xcut29 
transform 1 0 1008 0 1 686
box 1008 686 1042 778
use SUNSAR_cut_M1M3_2x1 xcut30 
transform 1 0 1222 0 1 1325
box 1222 1325 1314 1359
use SUNSAR_cut_M2M3_1x2 xcut31 
transform 1 0 1008 0 1 1298
box 1008 1298 1042 1390
use SUNSAR_cut_M1M3_2x1 xcut32 
transform 1 0 1222 0 1 1019
box 1222 1019 1314 1053
use SUNSAR_cut_M2M3_1x2 xcut33 
transform 1 0 1008 0 1 992
box 1008 992 1042 1084
use SUNSAR_cut_M1M3_2x1 xcut34 
transform 1 0 1222 0 1 407
box 1222 407 1314 441
use SUNSAR_cut_M2M3_1x2 xcut35 
transform 1 0 1008 0 1 380
box 1008 380 1042 472
use SUNSAR_cut_M1M3_2x1 xcut36 
transform 1 0 1222 0 1 7045
box 1222 7045 1314 7079
use SUNSAR_cut_M2M3_1x2 xcut37 
transform 1 0 1008 0 1 7018
box 1008 7018 1042 7110
use SUNSAR_cut_M1M3_2x1 xcut38 
transform 1 0 1222 0 1 8575
box 1222 8575 1314 8609
use SUNSAR_cut_M2M3_1x2 xcut39 
transform 1 0 1008 0 1 8548
box 1008 8548 1042 8640
use SUNSAR_cut_M1M3_2x1 xcut40 
transform 1 0 1222 0 1 7657
box 1222 7657 1314 7691
use SUNSAR_cut_M2M3_1x2 xcut41 
transform 1 0 1008 0 1 7630
box 1008 7630 1042 7722
use SUNSAR_cut_M1M3_2x1 xcut42 
transform 1 0 1222 0 1 8269
box 1222 8269 1314 8303
use SUNSAR_cut_M2M3_1x2 xcut43 
transform 1 0 1008 0 1 8242
box 1008 8242 1042 8334
use SUNSAR_cut_M1M3_2x1 xcut44 
transform 1 0 1222 0 1 7963
box 1222 7963 1314 7997
use SUNSAR_cut_M2M3_1x2 xcut45 
transform 1 0 1008 0 1 7936
box 1008 7936 1042 8028
use SUNSAR_cut_M1M3_2x1 xcut46 
transform 1 0 1222 0 1 7351
box 1222 7351 1314 7385
use SUNSAR_cut_M2M3_1x2 xcut47 
transform 1 0 1008 0 1 7324
box 1008 7324 1042 7416
use SUNSAR_cut_M1M3_2x1 xcut48 
transform 1 0 1222 0 1 10517
box 1222 10517 1314 10551
use SUNSAR_cut_M2M3_1x2 xcut49 
transform 1 0 914 0 1 10490
box 914 10490 948 10582
use SUNSAR_cut_M1M3_2x1 xcut50 
transform 1 0 1222 0 1 12047
box 1222 12047 1314 12081
use SUNSAR_cut_M2M3_1x2 xcut51 
transform 1 0 914 0 1 12020
box 914 12020 948 12112
use SUNSAR_cut_M1M3_2x1 xcut52 
transform 1 0 1222 0 1 11129
box 1222 11129 1314 11163
use SUNSAR_cut_M2M3_1x2 xcut53 
transform 1 0 914 0 1 11102
box 914 11102 948 11194
use SUNSAR_cut_M1M3_2x1 xcut54 
transform 1 0 1222 0 1 11741
box 1222 11741 1314 11775
use SUNSAR_cut_M2M3_1x2 xcut55 
transform 1 0 914 0 1 11714
box 914 11714 948 11806
use SUNSAR_cut_M1M3_2x1 xcut56 
transform 1 0 1222 0 1 11435
box 1222 11435 1314 11469
use SUNSAR_cut_M2M3_1x2 xcut57 
transform 1 0 914 0 1 11408
box 914 11408 948 11500
use SUNSAR_cut_M1M3_2x1 xcut58 
transform 1 0 1222 0 1 10823
box 1222 10823 1314 10857
use SUNSAR_cut_M2M3_1x2 xcut59 
transform 1 0 914 0 1 10796
box 914 10796 948 10888
use SUNSAR_cut_M1M3_2x1 xcut60 
transform 1 0 1222 0 1 1837
box 1222 1837 1314 1871
use SUNSAR_cut_M2M3_1x2 xcut61 
transform 1 0 820 0 1 1810
box 820 1810 854 1902
use SUNSAR_cut_M1M3_2x1 xcut62 
transform 1 0 1222 0 1 3367
box 1222 3367 1314 3401
use SUNSAR_cut_M2M3_1x2 xcut63 
transform 1 0 820 0 1 3340
box 820 3340 854 3432
use SUNSAR_cut_M1M3_2x1 xcut64 
transform 1 0 1222 0 1 2449
box 1222 2449 1314 2483
use SUNSAR_cut_M2M3_1x2 xcut65 
transform 1 0 820 0 1 2422
box 820 2422 854 2514
use SUNSAR_cut_M1M3_2x1 xcut66 
transform 1 0 1222 0 1 3061
box 1222 3061 1314 3095
use SUNSAR_cut_M2M3_1x2 xcut67 
transform 1 0 820 0 1 3034
box 820 3034 854 3126
use SUNSAR_cut_M1M3_2x1 xcut68 
transform 1 0 1222 0 1 2755
box 1222 2755 1314 2789
use SUNSAR_cut_M2M3_1x2 xcut69 
transform 1 0 820 0 1 2728
box 820 2728 854 2820
use SUNSAR_cut_M1M3_2x1 xcut70 
transform 1 0 1222 0 1 2143
box 1222 2143 1314 2177
use SUNSAR_cut_M2M3_1x2 xcut71 
transform 1 0 820 0 1 2116
box 820 2116 854 2208
use SUNSAR_cut_M1M3_2x1 xcut72 
transform 1 0 1222 0 1 3879
box 1222 3879 1314 3913
use SUNSAR_cut_M2M3_1x2 xcut73 
transform 1 0 726 0 1 3852
box 726 3852 760 3944
use SUNSAR_cut_M1M3_2x1 xcut74 
transform 1 0 1222 0 1 9087
box 1222 9087 1314 9121
use SUNSAR_cut_M2M3_1x2 xcut75 
transform 1 0 632 0 1 9060
box 632 9060 666 9152
use SUNSAR_cut_M1M3_2x1 xcut76 
transform 1 0 1222 0 1 8781
box 1222 8781 1314 8815
use SUNSAR_cut_M2M3_1x2 xcut77 
transform 1 0 538 0 1 8754
box 538 8754 572 8846
use SUNSAR_cut_M1M3_2x1 xcut78 
transform 1 0 1222 0 1 10311
box 1222 10311 1314 10345
use SUNSAR_cut_M2M3_1x2 xcut79 
transform 1 0 538 0 1 10284
box 538 10284 572 10376
use SUNSAR_cut_M1M3_2x1 xcut80 
transform 1 0 1222 0 1 9393
box 1222 9393 1314 9427
use SUNSAR_cut_M2M3_1x2 xcut81 
transform 1 0 538 0 1 9366
box 538 9366 572 9458
use SUNSAR_cut_M1M3_2x1 xcut82 
transform 1 0 1222 0 1 10005
box 1222 10005 1314 10039
use SUNSAR_cut_M2M3_1x2 xcut83 
transform 1 0 538 0 1 9978
box 538 9978 572 10070
use SUNSAR_cut_M1M3_2x1 xcut84 
transform 1 0 1222 0 1 9699
box 1222 9699 1314 9733
use SUNSAR_cut_M2M3_1x2 xcut85 
transform 1 0 444 0 1 9672
box 444 9672 478 9764
use SUNSAR_cut_M1M3_2x1 xcut86 
transform 1 0 1222 0 1 4491
box 1222 4491 1314 4525
use SUNSAR_cut_M2M3_1x2 xcut87 
transform 1 0 350 0 1 4464
box 350 4464 384 4556
use SUNSAR_cut_M1M3_2x1 xcut88 
transform 1 0 1222 0 1 4797
box 1222 4797 1314 4831
use SUNSAR_cut_M2M3_1x2 xcut89 
transform 1 0 256 0 1 4770
box 256 4770 290 4862
use SUNSAR_cut_M1M3_2x1 xcut90 
transform 1 0 1222 0 1 4185
box 1222 4185 1314 4219
use SUNSAR_cut_M2M3_1x2 xcut91 
transform 1 0 162 0 1 4158
box 162 4158 196 4250
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 1222 0 1 5103
box 1222 5103 1314 5137
use SUNSAR_cut_M2M3_1x2 xcut93 
transform 1 0 68 0 1 5076
box 68 5076 102 5168
<< labels >>
flabel m1 s 1102 5282 1136 13888 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew signal bidirectional
flabel m1 s 1008 74 1042 13888 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew signal bidirectional
flabel m1 s 914 10490 948 13888 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew signal bidirectional
flabel m1 s 820 1810 854 13888 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew signal bidirectional
flabel m1 s 726 3852 760 13888 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew signal bidirectional
flabel m1 s 632 9060 666 13888 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew signal bidirectional
flabel m1 s 538 8754 572 13888 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew signal bidirectional
flabel m1 s 444 9672 478 13888 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew signal bidirectional
flabel m1 s 350 4464 384 13888 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew signal bidirectional
flabel m1 s 256 4770 290 13888 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew signal bidirectional
flabel m1 s 162 4158 196 13888 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew signal bidirectional
flabel m1 s 68 5076 102 13888 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew signal bidirectional
flabel m1 s 1386 0 5936 38 0 FreeSans 400 0 0 0 AVSS
port 14 nsew signal bidirectional
flabel m3 s 1386 12152 1424 13922 0 FreeSans 400 0 0 0 CTOP
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 68 0 5974 13922
<< end >>
