magic
tech sky130B
magscale 1 2
timestamp 1708383600
<< checkpaint >>
rect 0 0 2520 1408
<< locali >>
rect 1622 582 1690 826
rect 1622 934 1690 1178
rect 864 230 1032 298
rect 864 582 1032 650
rect 864 758 1032 826
rect 1032 230 1100 826
rect 1420 406 1656 474
rect 864 1286 1420 1354
rect 1420 406 1488 1354
rect 1656 54 1824 122
rect 1824 1198 2088 1266
rect 1824 54 1892 1266
rect 756 54 1764 122
rect 2412 132 2628 220
rect -108 132 108 220
rect 324 846 540 914
rect 324 494 540 562
rect 1980 142 2196 210
rect 324 142 540 210
rect 1548 406 1764 474
<< poly >>
rect 324 510 2196 546
rect 324 862 2196 898
rect 324 1214 2196 1250
<< m3 >>
rect 1548 0 1732 1408
rect 756 0 940 1408
rect 1548 0 1732 1408
rect 756 0 940 1408
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNSAR_NCHDL MN3 
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNSAR_PCHDL MP0 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_PCHDL MP2 
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNSAR_PCHDL MP3 
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 230
box 1548 230 1732 298
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 1548 0 1 1286
box 1548 1286 1732 1354
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 756 0 1 406
box 756 406 940 474
use SUNSAR_cut_M1M4_2x1 xcut3 
transform 1 0 756 0 1 934
box 756 934 940 1002
use SUNSAR_cut_M1M4_2x1 xcut4 
transform 1 0 756 0 1 1110
box 756 1110 940 1178
<< labels >>
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel locali s 324 846 540 914 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 324 494 540 562 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 1980 142 2196 210 0 FreeSans 400 0 0 0 RST_N
port 5 nsew signal bidirectional
flabel locali s 324 142 540 210 0 FreeSans 400 0 0 0 EN
port 3 nsew signal bidirectional
flabel locali s 1548 406 1764 474 0 FreeSans 400 0 0 0 ENO
port 4 nsew signal bidirectional
flabel m3 s 1548 0 1732 1408 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 756 0 940 1408 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 2520 0 1408
<< end >>
