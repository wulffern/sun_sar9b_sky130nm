magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 1260 440
<< locali >>
rect 432 115 516 149
rect 432 291 516 325
rect 516 115 828 149
rect 516 291 828 325
rect 516 115 550 325
rect 199 71 233 369
rect 1027 71 1061 369
rect 162 71 270 105
rect 378 115 486 149
rect 1206 66 1314 110
rect -54 66 54 110
<< poly >>
rect 162 79 1098 97
rect 162 167 1098 185
rect 162 255 1098 273
rect 162 343 1098 361
<< m3 >>
rect 774 0 874 440
rect 378 0 478 440
rect 774 0 874 440
rect 378 0 478 440
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 88
box 0 88 630 264
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 176
box 0 176 630 352
use SUNSAR_NCHDL MN3 
transform 1 0 0 0 1 264
box 0 264 630 440
use SUNSAR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNSAR_PCHDL MP1 
transform 1 0 630 0 1 88
box 630 88 1260 264
use SUNSAR_PCHDL MP2 
transform 1 0 630 0 1 176
box 630 176 1260 352
use SUNSAR_PCHDL MP3 
transform 1 0 630 0 1 264
box 630 264 1260 440
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 27
box 774 27 874 65
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 203
box 774 203 874 241
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 774 0 1 203
box 774 203 874 241
use SUNSAR_cut_M1M4_2x1 xcut3 
transform 1 0 774 0 1 379
box 774 379 874 417
use SUNSAR_cut_M1M4_2x1 xcut4 
transform 1 0 378 0 1 27
box 378 27 478 65
use SUNSAR_cut_M1M4_2x1 xcut5 
transform 1 0 378 0 1 203
box 378 203 478 241
use SUNSAR_cut_M1M4_2x1 xcut6 
transform 1 0 378 0 1 203
box 378 203 478 241
use SUNSAR_cut_M1M4_2x1 xcut7 
transform 1 0 378 0 1 379
box 378 379 478 417
<< labels >>
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 378 115 486 149 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 3 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 4 nsew signal bidirectional
flabel m3 s 774 0 874 440 0 FreeSans 400 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel m3 s 378 0 478 440 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 440
<< end >>
