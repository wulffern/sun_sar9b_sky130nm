* NGSPICE file created from SUNSAR_SAR9B_CV.ext - technology: sky130A

.subckt SUNSAR_RM1 A B 0
R0 A B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
.ends

.subckt SUNSAR_CAP32C_CV C1A C1B C2 C4 C8 C16 CTOP XRES1A/B 0 XRES1B/B AVSS
XXRES16 C16 XRES16/B 0 SUNSAR_RM1
XXRES2 C2 XRES2/B 0 SUNSAR_RM1
XXRES1A C1A XRES1A/B 0 SUNSAR_RM1
XXRES1B C1B XRES1B/B 0 SUNSAR_RM1
XXRES4 C4 XRES4/B 0 SUNSAR_RM1
XXRES8 C8 XRES8/B 0 SUNSAR_RM1
C0 XRES1A/B CTOP 3.637777f
C1 XRES2/B CTOP 7.010892f
C2 AVSS XRES16/B 10.460171f
C3 XRES8/B XRES16/B 0.1057f
C4 XRES8/B AVSS 7.113892f
C5 XRES4/B XRES16/B 0.063821f
C6 XRES4/B AVSS 5.459597f
C7 XRES1B/B XRES16/B 0.05157f
C8 XRES4/B XRES8/B 0.477132f
C9 XRES1B/B AVSS 4.270325f
C10 XRES16/B CTOP 55.2954f
C11 AVSS CTOP 11.093214f
C12 XRES1A/B XRES16/B 0.467299f
C13 XRES1A/B AVSS 4.264343f
C14 XRES2/B XRES16/B 0.470901f
C15 XRES8/B CTOP 27.705545f
C16 XRES2/B AVSS 4.595231f
C17 XRES1B/B XRES4/B 0.430616f
C18 XRES2/B XRES8/B 0.446669f
C19 XRES4/B CTOP 13.930625f
C20 XRES1B/B CTOP 3.637325f
C21 CTOP 0 7.97522f
C22 XRES16/B 0 4.882493f
C23 AVSS 0 16.502905f
C24 XRES8/B 0 4.160811f
C25 C8 0 0.111021f
C26 XRES4/B 0 3.74557f
C27 C4 0 0.111021f
C28 XRES1B/B 0 3.31589f
C29 C1B 0 0.12719f
C30 XRES1A/B 0 1.751233f
C31 C1A 0 0.12719f
C32 XRES2/B 0 3.488749f
C33 C2 0 0.111021f
C34 C16 0 0.111021f
.ends

.subckt SUNSAR_CDAC8_CV CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1>
+ CP<0> CTOP XC1/XRES1A/B CP<11> 0 AVSS
XXC128b<2> CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP XC128b<2>/XRES1A/B 0 XC128b<2>/XRES1B/B
+ AVSS SUNSAR_CAP32C_CV
XX16ab CP<5> CP<5> CP<5> CP<5> CP<4> CP<6> CTOP X16ab/XRES1A/B 0 X16ab/XRES1B/B AVSS
+ SUNSAR_CAP32C_CV
XXC64a<0> CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CTOP XC64a<0>/XRES1A/B 0 XC64a<0>/XRES1B/B
+ AVSS SUNSAR_CAP32C_CV
XXC0 CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP XC0/XRES1A/B 0 XC0/XRES1B/B AVSS
+ SUNSAR_CAP32C_CV
XXC1 CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP XC1/XRES1A/B 0 XC1/XRES1B/B AVSS
+ SUNSAR_CAP32C_CV
XXC64b<1> CP<9> CP<9> CP<9> CP<9> CP<9> CP<9> CTOP XC64b<1>/XRES1A/B 0 XC64b<1>/XRES1B/B
+ AVSS SUNSAR_CAP32C_CV
XXC128a<1> CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP XC128a<1>/XRES1A/B 0 XC128a<1>/XRES1B/B
+ AVSS SUNSAR_CAP32C_CV
XXC32a<0> AVSS CP<0> CP<1> CP<2> CP<3> CP<7> CTOP XC32a<0>/XRES1A/B 0 XC32a<0>/XRES1B/B
+ AVSS SUNSAR_CAP32C_CV
C0 XC64b<1>/XRES1B/B AVSS 0.094089f
C1 XC64b<1>/XRES1A/B X16ab/XRES1B/B 0.628951f
C2 CP<3> CP<4> 2.189413f
C3 CP<11> CP<5> 0.395544f
C4 CP<11> CP<6> 0.1009f
C5 CP<10> AVSS 0.759823f
C6 AVSS XC32a<0>/XRES1B/B 0.094089f
C7 CP<10> CP<7> 0.103863f
C8 CP<0> CP<1> 4.6508f
C9 XC64b<1>/XRES1A/B AVSS 0.094956f
C10 AVSS CTOP -4.036157f
C11 CP<0> CP<3> 0.089475f
C12 CP<0> CP<2> 0.276335f
C13 CP<9> AVSS 0.097224f
C14 AVSS XC128a<1>/XRES1B/B 0.094089f
C15 XC128b<2>/XRES1A/B XC128a<1>/XRES1B/B 0.628951f
C16 CP<6> CP<5> 3.024884f
C17 CP<7> CP<4> 0.082973f
C18 CP<10> CP<8> 2.855174f
C19 AVSS XC128a<1>/XRES1A/B 0.094956f
C20 CP<3> CP<5> 0.232224f
C21 CP<8> CTOP 0.112463f
C22 CP<11> AVSS 1.417505f
C23 CP<7> CP<0> 0.089189f
C24 CP<3> CP<1> 0.253055f
C25 CP<2> CP<1> 4.734883f
C26 XC1/XRES1B/B AVSS 0.094089f
C27 CP<9> CP<8> 1.80154f
C28 CP<2> CP<3> 4.987515f
C29 CP<8> CP<4> 0.086534f
C30 AVSS CP<5> 0.064356f
C31 CP<7> CP<5> 0.415707f
C32 XC0/XRES1A/B AVSS 0.094956f
C33 CP<7> CP<6> 2.585879f
C34 CP<10> CTOP 0.236926f
C35 CP<0> CP<8> 0.087696f
C36 CP<7> CP<1> 0.225261f
C37 CP<9> CP<10> 2.280731f
C38 CP<7> CP<3> 0.602343f
C39 AVSS XC32a<0>/XRES1A/B 0.094956f
C40 CP<7> CP<2> 0.087928f
C41 CP<9> CTOP 0.073803f
C42 CP<10> CP<4> 0.086632f
C43 XC64a<0>/XRES1A/B XC1/XRES1B/B 0.62895f
C44 CP<8> CP<5> 0.349544f
C45 XC128b<2>/XRES1B/B AVSS 0.094089f
C46 X16ab/XRES1B/B AVSS 0.094089f
C47 XC128a<1>/XRES1A/B XC32a<0>/XRES1B/B 0.62895f
C48 XC128b<2>/XRES1B/B X16ab/XRES1A/B 0.62895f
C49 CP<8> CP<6> 0.087273f
C50 CP<10> CP<0> 0.099397f
C51 CP<10> CP<11> 5.253161f
C52 CP<8> CP<1> 0.08638f
C53 CP<8> CP<3> 0.086451f
C54 XC128b<2>/XRES1A/B AVSS 0.094956f
C55 X16ab/XRES1A/B AVSS 0.094956f
C56 CP<8> CP<2> 0.086407f
C57 CP<11> CTOP 0.226487f
C58 XC64a<0>/XRES1B/B XC32a<0>/XRES1A/B 0.628951f
C59 XC64b<1>/XRES1B/B XC0/XRES1A/B 0.62895f
C60 CP<9> CP<11> 0.702233f
C61 CP<10> CP<5> 0.461689f
C62 CP<10> CP<6> 0.08676f
C63 CP<11> CP<4> 0.100006f
C64 CP<10> CP<1> 0.098065f
C65 CP<10> CP<3> 0.098862f
C66 CP<8> AVSS 0.141321f
C67 XC64a<0>/XRES1B/B AVSS 0.094089f
C68 CP<10> CP<2> 0.098672f
C69 CP<9> CP<5> 0.144727f
C70 CP<7> CP<8> 5.335522f
C71 CP<11> CP<0> 0.094714f
C72 CP<5> CP<4> 2.571549f
C73 CP<6> CP<4> 0.08351f
C74 XC64a<0>/XRES1A/B AVSS 0.094956f
C75 CP<10> 0 7.076044f
C76 CP<8> 0 4.111091f
C77 CP<7> 0 0.984698f
C78 CP<1> 0 1.553364f
C79 CP<3> 0 1.105384f
C80 CP<2> 0 0.987259f
C81 CP<0> 0 1.541327f
C82 CP<11> 0 5.570052f
C83 CP<5> 0 2.62574f
C84 CP<6> 0 0.780529f
C85 CP<4> 0 0.889614f
C86 CP<9> 0 2.620203f
C87 XC32a<0>/XRES16/B 0 4.882493f
C88 XC32a<0>/XRES8/B 0 4.160811f
C89 XC32a<0>/XRES4/B 0 3.74557f
C90 XC32a<0>/XRES1B/B 0 3.31589f
C91 XC32a<0>/XRES1A/B 0 1.751233f
C92 XC32a<0>/XRES2/B 0 3.488749f
C93 XC128a<1>/XRES16/B 0 4.882493f
C94 XC128a<1>/XRES8/B 0 4.160811f
C95 XC128a<1>/XRES4/B 0 3.74557f
C96 XC128a<1>/XRES1B/B 0 3.31589f
C97 XC128a<1>/XRES1A/B 0 1.751233f
C98 XC128a<1>/XRES2/B 0 3.488749f
C99 XC64b<1>/XRES16/B 0 4.882493f
C100 XC64b<1>/XRES8/B 0 4.160811f
C101 XC64b<1>/XRES4/B 0 3.74557f
C102 XC64b<1>/XRES1B/B 0 3.31589f
C103 XC64b<1>/XRES1A/B 0 1.751233f
C104 XC64b<1>/XRES2/B 0 3.488749f
C105 CTOP 0 37.11138f
C106 XC1/XRES16/B 0 4.882493f
C107 AVSS 0 0.100432p
C108 XC1/XRES8/B 0 4.160811f
C109 XC1/XRES4/B 0 3.74557f
C110 XC1/XRES1B/B 0 3.31589f
C111 XC1/XRES1A/B 0 1.751233f
C112 XC1/XRES2/B 0 3.488749f
C113 XC0/XRES16/B 0 4.882493f
C114 XC0/XRES8/B 0 4.160811f
C115 XC0/XRES4/B 0 3.74557f
C116 XC0/XRES1B/B 0 3.31589f
C117 XC0/XRES1A/B 0 1.751233f
C118 XC0/XRES2/B 0 3.488749f
C119 XC64a<0>/XRES16/B 0 4.882493f
C120 XC64a<0>/XRES8/B 0 4.160811f
C121 XC64a<0>/XRES4/B 0 3.74557f
C122 XC64a<0>/XRES1B/B 0 3.31589f
C123 XC64a<0>/XRES1A/B 0 1.751233f
C124 XC64a<0>/XRES2/B 0 3.488749f
C125 X16ab/XRES16/B 0 4.882493f
C126 X16ab/XRES8/B 0 4.160811f
C127 X16ab/XRES4/B 0 3.74557f
C128 X16ab/XRES1B/B 0 3.31589f
C129 X16ab/XRES1A/B 0 1.751233f
C130 X16ab/XRES2/B 0 3.488749f
C131 XC128b<2>/XRES16/B 0 4.882493f
C132 XC128b<2>/XRES8/B 0 4.160811f
C133 XC128b<2>/XRES4/B 0 3.74557f
C134 XC128b<2>/XRES1B/B 0 3.31589f
C135 XC128b<2>/XRES1A/B 0 1.751233f
C136 XC128b<2>/XRES2/B 0 3.488749f
.ends

.subckt SUNSAR_PCHDL D G S B 0 a_216_n18# a_216_334#
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 a_216_n18# B 0.330729f
C1 a_216_334# B 0.331144f
C2 D S 0.050207f
C3 G B 0.341895f
C4 a_216_n18# G 0.067588f
C5 G a_216_334# 0.066018f
C6 G 0 0.073301f
C7 B 0 2.80584f
C8 a_216_n18# 0 0.091271f
C9 a_216_334# 0 0.091271f
.ends

.subckt SUNSAR_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 G a_324_n18# 0.066018f
C1 S D 0.050207f
C2 G a_324_334# 0.067588f
C3 S B 0.06638f
C4 G B 0.415197f
C5 D B 0.06638f
C6 a_324_n18# B 0.422415f
C7 a_324_334# B 0.422f
.ends

.subckt SUNSAR_NDX1_CV Y AVDD AVSS MN1/a_324_334# B A BULKP BULKN MP0/a_216_n18# MP1/a_216_334#
+ MN0/a_324_n18#
XMP0 Y A AVDD BULKP BULKN MP0/a_216_n18# B SUNSAR_PCHDL
XMP1 AVDD B Y BULKP BULKN A MP1/a_216_334# SUNSAR_PCHDL
XMN0 MN1/S A AVSS BULKN MN0/a_324_n18# B SUNSAR_NCHDL
XMN1 Y B MN1/S BULKN A MN1/a_324_334# SUNSAR_NCHDL
C0 Y AVDD 0.078555f
C1 BULKP AVDD 0.15616f
C2 A BULKP -0.246413f
C3 Y B 0.059989f
C4 AVDD AVSS 0.072347f
C5 B BULKP -0.247362f
C6 AVSS BULKN 0.399663f
C7 MN1/a_324_334# BULKN 0.422f
C8 AVDD BULKN 0.333494f
C9 MN0/a_324_n18# BULKN 0.422415f
C10 Y BULKN 0.252959f
C11 B BULKN 0.538314f
C12 BULKP BULKN 3.595964f
C13 A BULKN 0.539194f
C14 MP1/a_216_334# BULKN 0.091338f
C15 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_NRX1_CV AVSS MN1/a_324_334# B BULKP BULKN MP0/a_216_n18# Y MP1/a_216_334#
+ AVDD A MN0/a_324_n18#
XMP0 MP1/S A AVDD BULKP BULKN MP0/a_216_n18# B SUNSAR_PCHDL
XMP1 Y B MP1/S BULKP BULKN A MP1/a_216_334# SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# B SUNSAR_NCHDL
XMN1 AVSS B Y BULKN A MN1/a_324_334# SUNSAR_NCHDL
C0 AVDD AVSS 0.072522f
C1 BULKP Y 0.076318f
C2 AVDD BULKP 0.12362f
C3 BULKP A -0.246413f
C4 B Y 0.059989f
C5 B BULKP -0.247362f
C6 AVSS Y 0.114122f
C7 Y BULKN 0.247181f
C8 MN1/a_324_334# BULKN 0.422f
C9 AVSS BULKN 0.513412f
C10 MN0/a_324_n18# BULKN 0.422415f
C11 AVDD BULKN 0.264177f
C12 B BULKN 0.538314f
C13 BULKP BULKN 3.595964f
C14 MP1/a_216_334# BULKN 0.091338f
C15 A BULKN 0.539194f
C16 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_IVX1_CV BULKP AVSS Y BULKN MP0/a_216_n18# MP0/a_216_334# AVDD A MN0/a_324_n18#
+ MN0/a_324_334#
XMP0 Y A AVDD BULKP BULKN MP0/a_216_n18# MP0/a_216_334# SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 Y BULKP 0.061437f
C1 AVDD BULKP 0.104456f
C2 A BULKP 0.109299f
C3 AVSS AVDD 0.0519f
C4 AVSS BULKN 0.374279f
C5 MN0/a_324_n18# BULKN 0.422415f
C6 MN0/a_324_334# BULKN 0.422f
C7 AVDD BULKN 0.252941f
C8 A BULKN 0.631634f
C9 Y BULKN 0.268384f
C10 BULKP BULKN 2.80697f
C11 MP0/a_216_n18# BULKN 0.091338f
C12 MP0/a_216_334# BULKN 0.091338f
.ends

.subckt SUNSAR_TAPCELLB_CV AVSS MN1/a_324_n18# MN1/a_324_334# MP1/a_216_334# MP1/a_216_n18#
+ AVDD
XMP1 AVDD AVDD AVDD AVDD AVSS MP1/a_216_n18# MP1/a_216_334# SUNSAR_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNSAR_NCHDL
C0 AVDD AVSS 0.105819f
C1 AVSS 0 1.05597f
C2 MN1/a_324_n18# 0 0.422415f
C3 MN1/a_324_334# 0 0.422f
C4 AVDD 0 3.141198f
C5 MP1/a_216_n18# 0 0.091271f
C6 MP1/a_216_334# 0 0.091271f
.ends

.subckt SUNSAR_SARKICKHX1_CV CI BULKP AVDD AVSS MP6_DMY/a_216_334# MN6/a_324_334#
+ MP0/S CKN MP0/a_216_n18# CK BULKN MN0/a_324_n18#
XMP1_DMY AVDD AVDD AVDD BULKP BULKN CKN AVDD SUNSAR_PCHDL
XMP4_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
XMP0 AVDD CKN MP0/S BULKP BULKN MP0/a_216_n18# AVDD SUNSAR_PCHDL
XMN0 MP0/S CKN AVSS BULKN MN0/a_324_n18# CI SUNSAR_NCHDL
XMN1 MP0/S CI MP0/S BULKN CKN CI SUNSAR_NCHDL
XMN2 MP0/S CI MP0/S BULKN CI CI SUNSAR_NCHDL
XMN3 MP0/S CI MP0/S BULKN CI CI SUNSAR_NCHDL
XMN4 MP0/S CI MP0/S BULKN CI CI SUNSAR_NCHDL
XMN6 AVDD CK MP0/S BULKN CI MN6/a_324_334# SUNSAR_NCHDL
XMN5 MP0/S CI MP0/S BULKN CI CK SUNSAR_NCHDL
XMP3_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
XMP6_DMY AVDD AVDD AVDD BULKP BULKN AVDD MP6_DMY/a_216_334# SUNSAR_PCHDL
XMP2_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
XMP5_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
C0 CKN MP0/S 0.058228f
C1 BULKP MP0/S 0.11694f
C2 AVDD MP0/S 0.103723f
C3 AVDD AVSS 0.185084f
C4 CKN BULKP -0.227092f
C5 AVDD BULKP -3.512327f
C6 MP0/S AVSS 0.214157f
C7 CI MP0/S -0.056784f
C8 CI AVSS 0.053147f
C9 BULKP BULKN 7.544365f
C10 MP6_DMY/a_216_334# BULKN 0.091338f
C11 AVDD BULKN 0.750023f
C12 CK BULKN 0.372036f
C13 MN6/a_324_334# BULKN 0.422f
C14 CI BULKN 1.791641f
C15 AVSS BULKN 0.562555f
C16 MN0/a_324_n18# BULKN 0.422415f
C17 MP0/S BULKN 0.370985f
C18 MP0/a_216_n18# BULKN 0.091338f
C19 CKN BULKN 0.56349f
.ends

.subckt SUNSAR_SARCMPHX1_CV CI CK VMR N2 AVDD AVSS MP6/a_216_334# MN6/a_324_334# BULKN
+ MP0/a_216_n18# BULKP CO MN0/a_324_n18# N1
XMP0 AVDD CK N1 BULKP BULKN MP0/a_216_n18# CK SUNSAR_PCHDL
XMP1 N2 CK AVDD BULKP BULKN CK AVDD SUNSAR_PCHDL
XMN0 N1 CK AVSS BULKN MN0/a_324_n18# CI SUNSAR_NCHDL
XMP2 AVDD AVDD N2 BULKP BULKN CK CK SUNSAR_PCHDL
XMN1 N2 CI N1 BULKN CK CI SUNSAR_NCHDL
XMP3 CO CK AVDD BULKP BULKN AVDD VMR SUNSAR_PCHDL
XMP4 AVDD VMR CO BULKP BULKN CK VMR SUNSAR_PCHDL
XMN2 N1 CI N2 BULKN CI CI SUNSAR_NCHDL
XMP5 CO VMR AVDD BULKP BULKN VMR VMR SUNSAR_PCHDL
XMN3 N2 CI N1 BULKN CI CI SUNSAR_NCHDL
XMN4 N1 CI N2 BULKN CI CI SUNSAR_NCHDL
XMP6 AVDD VMR CO BULKP BULKN VMR MP6/a_216_334# SUNSAR_PCHDL
XMN5 N2 CI N1 BULKN CI VMR SUNSAR_NCHDL
XMN6 CO VMR N2 BULKN CI MN6/a_324_334# SUNSAR_NCHDL
C0 N1 CI 0.175052f
C1 N2 CO 0.076147f
C2 BULKP CK -1.349649f
C3 BULKP CO 0.063159f
C4 N2 AVSS 0.099131f
C5 CO VMR 0.076819f
C6 AVDD CK 0.064755f
C7 AVDD CO 0.223072f
C8 BULKP N2 0.063625f
C9 AVDD AVSS 0.161411f
C10 N1 CK 0.072917f
C11 N1 AVSS 0.16219f
C12 BULKP VMR -1.552184f
C13 AVDD N2 0.080291f
C14 CI AVSS 0.05721f
C15 AVDD BULKP -0.437744f
C16 N1 N2 0.189549f
C17 AVDD VMR 0.051752f
C18 N1 BULKP 0.069686f
C19 N1 AVDD 0.058844f
C20 AVSS BULKN 0.540993f
C21 MN6/a_324_334# BULKN 0.422f
C22 VMR BULKN 0.606867f
C23 MP6/a_216_334# BULKN 0.091338f
C24 CI BULKN 1.771056f
C25 CK BULKN 0.626869f
C26 CO BULKN 0.213838f
C27 N2 BULKN 0.221339f
C28 BULKP BULKN 7.544966f
C29 MN0/a_324_n18# BULKN 0.422415f
C30 AVDD BULKN 0.618349f
C31 N1 BULKN 0.369132f
C32 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_IVX4_CV AVDD AVSS MP3/a_216_334# MN3/a_324_334# BULKN BULKP MP0/a_216_n18#
+ Y A MN0/a_324_n18#
XMP0 Y A AVDD BULKP BULKN MP0/a_216_n18# A SUNSAR_PCHDL
XMP1 AVDD A Y BULKP BULKN A A SUNSAR_PCHDL
XMP2 Y A AVDD BULKP BULKN A A SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# A SUNSAR_NCHDL
XMP3 AVDD A Y BULKP BULKN A MP3/a_216_334# SUNSAR_PCHDL
XMN1 AVSS A Y BULKN A A SUNSAR_NCHDL
XMN2 Y A AVSS BULKN A A SUNSAR_NCHDL
XMN3 AVSS A Y BULKN A MN3/a_324_334# SUNSAR_NCHDL
C0 Y A 0.147008f
C1 AVDD Y 0.147387f
C2 Y AVSS 0.177209f
C3 AVDD A 0.065686f
C4 AVSS A 0.065557f
C5 BULKP A -1.606473f
C6 AVDD AVSS 0.133497f
C7 BULKP AVDD 0.168357f
C8 A BULKN 2.062361f
C9 AVSS BULKN 0.629948f
C10 MN3/a_324_334# BULKN 0.422f
C11 MP3/a_216_334# BULKN 0.091338f
C12 Y BULKN 0.278637f
C13 MN0/a_324_n18# BULKN 0.422415f
C14 AVDD BULKN 0.379723f
C15 BULKP BULKN 5.176431f
C16 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARCMPX1_CV CPI CNI CK_CMP XA12/Y XA3/CO XA3a/A CK_SAMPLE XA9/A CPO
+ DONE AVSS CNO AVDD
XXA10 XA9/A AVDD AVSS XA11/MN0/a_324_n18# XA12/Y XA11/Y AVDD AVSS XA9/MP0/a_216_334#
+ XA11/MP0/a_216_n18# XA9/MN0/a_324_334# SUNSAR_NDX1_CV
XXA11 AVSS XA12/MN0/a_324_n18# DONE AVDD AVSS XA11/MP0/a_216_n18# XA11/Y XA12/MP0/a_216_n18#
+ AVDD CK_SAMPLE XA11/MN0/a_324_n18# SUNSAR_NRX1_CV
XXA12 AVDD AVSS XA12/Y AVSS XA12/MP0/a_216_n18# XA13/MP1/a_216_n18# AVDD CK_CMP XA12/MN0/a_324_n18#
+ XA13/MN1/a_324_n18# SUNSAR_IVX1_CV
XXA13 AVSS XA13/MN1/a_324_n18# XA13/MN1/a_324_334# XA13/MP1/a_216_334# XA13/MP1/a_216_n18#
+ AVDD SUNSAR_TAPCELLB_CV
XXA0 AVSS XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ AVDD SUNSAR_TAPCELLB_CV
XXA1 CPI AVDD AVDD AVSS XA2/MP0/a_216_n18# XA2/MN0/a_324_n18# XA1/MP0/S XA9/A XA1/MP0/a_216_n18#
+ XA9/Y AVSS XA1/MN0/a_324_n18# SUNSAR_SARKICKHX1_CV
XXA2 CPI XA9/Y XA3/CO XA2/N2 AVDD AVSS XA2/MP6/a_216_334# XA2/MN6/a_324_334# AVSS
+ XA2/MP0/a_216_n18# AVDD XA3a/A XA2/MN0/a_324_n18# XA3/N1 SUNSAR_SARCMPHX1_CV
XXA3 CNI XA9/Y XA3a/A XA3/N2 AVDD AVSS XA4/MP0/a_216_n18# XA4/MN0/a_324_n18# AVSS
+ XA3/MP0/a_216_n18# AVDD XA3/CO XA3/MN0/a_324_n18# XA3/N1 SUNSAR_SARCMPHX1_CV
XXA4 CNI AVDD AVDD AVSS XA9/MP0/a_216_n18# XA9/MN0/a_324_n18# XA4/MP0/S XA9/A XA4/MP0/a_216_n18#
+ XA9/Y AVSS XA4/MN0/a_324_n18# SUNSAR_SARKICKHX1_CV
XXA3a AVDD AVSS XA3/MP0/a_216_n18# XA3/MN0/a_324_n18# AVSS AVDD XA3a/MP0/a_216_n18#
+ CNO XA3a/A XA3a/MN0/a_324_n18# SUNSAR_IVX4_CV
XXA2a AVDD AVSS XA3a/MP0/a_216_n18# XA3a/MN0/a_324_n18# AVSS AVDD XA2/MP6/a_216_334#
+ CPO XA3/CO XA2/MN6/a_324_334# SUNSAR_IVX4_CV
XXA9 AVDD AVSS XA9/Y AVSS XA9/MP0/a_216_n18# XA9/MP0/a_216_334# AVDD XA9/A XA9/MN0/a_324_n18#
+ XA9/MN0/a_324_334# SUNSAR_IVX1_CV
C0 XA12/Y AVDD 0.491363f
C1 XA9/Y CNI 0.382485f
C2 XA11/Y AVDD 0.055398f
C3 XA2/MP0/a_216_n18# AVDD -0.312114f
C4 XA11/Y XA9/A 0.268591f
C5 XA9/Y XA3/CO 0.24121f
C6 XA9/MP0/a_216_334# AVDD -0.311437f
C7 XA1/MP0/S AVDD 0.073206f
C8 XA3a/A XA3/CO 1.092423f
C9 XA3/N1 AVDD 0.19591f
C10 XA1/MP0/a_216_n18# AVDD -0.312114f
C11 XA3/N1 CNO 0.113873f
C12 XA2/MP6/a_216_334# AVDD -0.313651f
C13 XA4/MP0/a_216_n18# AVDD -0.312115f
C14 AVDD XA9/MP0/a_216_n18# -0.312114f
C15 XA3/N1 CPO 0.068565f
C16 CPI XA9/Y 0.27081f
C17 XA9/A AVDD 0.190387f
C18 XA9/Y XA3a/A 0.391167f
C19 AVDD XA3/MP0/a_216_n18# -0.313502f
C20 XA12/Y CK_SAMPLE 0.106092f
C21 CK_CMP DONE 0.058881f
C22 XA11/Y CK_SAMPLE 0.050093f
C23 XA3/N1 XA3/CO 0.289212f
C24 XA9/A CNI 0.362147f
C25 AVDD XA3/CO 1.186392f
C26 XA12/Y CK_CMP 0.05138f
C27 XA4/MP0/S XA3/CO 0.095491f
C28 XA9/A XA3/CO 0.141462f
C29 XA11/Y XA12/Y 0.130476f
C30 XA3/N1 XA9/Y 0.106124f
C31 XA3/N1 CPI 0.115376f
C32 XA9/Y AVDD 0.164538f
C33 XA3/N1 XA3a/A 0.309118f
C34 XA9/A XA9/Y 1.524979f
C35 AVDD XA3a/MP0/a_216_n18# -0.312395f
C36 XA9/A CPI 0.297822f
C37 AVDD XA3a/A 0.915439f
C38 XA12/MP0/a_216_n18# AVDD -0.312932f
C39 XA11/MP0/a_216_n18# AVDD -0.313072f
C40 XA9/A XA3a/A 0.136678f
C41 XA13/MP1/a_216_n18# AVDD -0.312114f
C42 XA3a/A CPO 0.108133f
C43 XA9/MN0/a_324_n18# AVSS 0.355024f
C44 XA3/CO AVSS 2.700815f
C45 CPO AVSS 0.178234f
C46 XA2/MN6/a_324_334# AVSS 0.353564f
C47 XA3a/A AVSS 2.52171f
C48 XA3/MN0/a_324_n18# AVSS 0.353564f
C49 CNO AVSS 0.179699f
C50 XA3a/MN0/a_324_n18# AVSS 0.353564f
C51 XA4/MN0/a_324_n18# AVSS 0.353572f
C52 XA4/MP0/S AVSS 0.414246f
C53 CNI AVSS 3.623488f
C54 XA3/N2 AVSS 0.246915f
C55 XA9/Y AVSS 4.611802f
C56 XA2/N2 AVSS 0.246915f
C57 XA2/MN0/a_324_n18# AVSS 0.353633f
C58 XA3/N1 AVSS 1.209705f
C59 AVDD AVSS 46.259968f
C60 CPI AVSS 3.747972f
C61 XA1/MN0/a_324_n18# AVSS 0.35614f
C62 XA1/MP0/S AVSS 0.422681f
C63 XA9/A AVSS 4.714037f
C64 XA0/MN1/a_324_n18# AVSS 0.422415f
C65 XA0/MP1/a_216_n18# AVSS 0.091271f
C66 XA13/MN1/a_324_334# AVSS 0.422f
C67 XA13/MP1/a_216_334# AVSS 0.091271f
C68 XA13/MN1/a_324_n18# AVSS 0.35614f
C69 CK_CMP AVSS 0.538443f
C70 XA12/MN0/a_324_n18# AVSS 0.356848f
C71 XA11/MN0/a_324_n18# AVSS 0.354112f
C72 DONE AVSS 0.474555f
C73 CK_SAMPLE AVSS 0.470113f
C74 XA9/MN0/a_324_334# AVSS 0.355615f
C75 XA12/Y AVSS 0.688598f
C76 XA11/Y AVSS 0.835691f
.ends

.subckt SUNSAR_NCHDLR D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 D S 0.050207f
C1 a_324_n18# G 0.066018f
C2 a_324_334# G 0.067588f
C3 S B 0.06638f
C4 G B 0.415197f
C5 D B 0.06638f
C6 a_324_n18# B 0.422415f
C7 a_324_334# B 0.422f
.ends

.subckt SUNSAR_CAP_BSSW_CV A B 0
R0 A m3_6948_120# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
R1 m3_252_280# B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
C0 A B 65.019196f
C1 m3_6948_120# B 0.172147f
C2 m3_6876_120# B 0.0666f
C3 m3_324_280# A 0.0666f
C4 m3_252_280# A 0.105547f
C5 B 0 13.2906f
C6 A 0 13.2887f
.ends

.subckt SUNSAR_CAP_BSSW5_CV B 0 A
XXCAPB0 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB1 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB2 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB3 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB4 A B 0 SUNSAR_CAP_BSSW_CV
C0 A B 54.00426f
C1 B 0 54.06679f
C2 A 0 55.079098f
.ends

.subckt SUNSAR_TIEH_CV Y BULKP AVDD AVSS BULKN MP0/a_216_n18# MP0/a_216_334# MP0/G
+ MN0/a_324_n18# MN0/a_324_334#
XMP0 Y MP0/G AVDD BULKP BULKN MP0/a_216_n18# MP0/a_216_334# SUNSAR_PCHDL
XMN0 MP0/G MP0/G AVSS BULKN MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.107492f
C1 BULKP MP0/G 0.112786f
C2 AVDD AVSS 0.0519f
C3 MP0/G AVSS 0.058774f
C4 AVSS BULKN 0.374633f
C5 MN0/a_324_n18# BULKN 0.422415f
C6 MN0/a_324_334# BULKN 0.422f
C7 AVDD BULKN 0.255369f
C8 MP0/G BULKN 0.790179f
C9 BULKP BULKN 2.806854f
C10 MP0/a_216_n18# BULKN 0.091338f
C11 MP0/a_216_334# BULKN 0.091338f
.ends

.subckt SUNSAR_TIEL_CV BULKP AVDD AVSS BULKN Y MP0/a_216_n18# MP0/a_216_334# MP0/G
+ MN0/a_324_n18# MN0/a_324_334#
XMP0 MP0/G MP0/G AVDD BULKP BULKN MP0/a_216_n18# MP0/a_216_334# SUNSAR_PCHDL
XMN0 Y MP0/G AVSS BULKN MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 MP0/G AVDD 0.05882f
C1 BULKP AVDD 0.104999f
C2 BULKP MP0/G 0.161174f
C3 AVDD AVSS 0.0519f
C4 AVSS BULKN 0.377294f
C5 Y BULKN 0.05974f
C6 MN0/a_324_n18# BULKN 0.422415f
C7 MN0/a_324_334# BULKN 0.422f
C8 AVDD BULKN 0.255397f
C9 MP0/G BULKN 0.708387f
C10 BULKP BULKN 2.806659f
C11 MP0/a_216_n18# BULKN 0.091338f
C12 MP0/a_216_334# BULKN 0.091338f
.ends

.subckt SUNSAR_TGPD_CV AVDD AVSS MP2/B MN2/a_324_334# MP0/S B MP0/a_216_n18# A 0 C
+ MP2/a_216_334# MN0/a_324_n18#
XMP1_DMY B AVDD AVDD MP2/B 0 C C SUNSAR_PCHDL
XMP0 AVDD C MP0/S MP2/B 0 MP0/a_216_n18# AVDD SUNSAR_PCHDL
XMP2 A C B MP2/B 0 AVDD MP2/a_216_334# SUNSAR_PCHDL
XMN0 AVSS C MP0/S 0 MN0/a_324_n18# C SUNSAR_NCHDL
XMN1 B C AVSS 0 C MP0/S SUNSAR_NCHDL
XMN2 A MP0/S B 0 C MN2/a_324_334# SUNSAR_NCHDL
C0 MP2/B C -0.388363f
C1 C AVDD 0.071397f
C2 AVSS AVDD 0.092101f
C3 MP2/B MP0/S 0.064367f
C4 MP0/S C 0.148714f
C5 B A 0.108f
C6 MP0/S AVSS 0.096157f
C7 MP0/S B 0.056087f
C8 MP2/B AVDD -0.503371f
C9 AVDD 0 0.485958f
C10 C 0 0.995572f
C11 AVSS 0 0.359707f
C12 A 0 0.204323f
C13 MN2/a_324_334# 0 0.422f
C14 B 0 0.060014f
C15 MP0/S 0 0.747699f
C16 MN0/a_324_n18# 0 0.422415f
C17 MP2/a_216_334# 0 0.091338f
C18 MP2/B 0 4.387254f
C19 MP0/a_216_n18# 0 0.091338f
.ends

.subckt SUNSAR_SARBSSWCTRL_CV GN GNG TIE_H AVDD AVSS MN1/a_324_334# C BULKP BULKN
+ MP0/a_216_n18# MP1/a_216_334# MN0/a_324_n18#
XMP0 GNG C GN BULKP BULKN MP0/a_216_n18# GN SUNSAR_PCHDL
XMP1 AVDD GN GNG BULKP BULKN C MP1/a_216_334# SUNSAR_PCHDL
XMN0 MN1/S C AVSS BULKN MN0/a_324_n18# TIE_H SUNSAR_NCHDL
XMN1 GN TIE_H MN1/S BULKN C MN1/a_324_334# SUNSAR_NCHDL
C0 AVDD AVSS 0.060449f
C1 GN AVSS 0.083748f
C2 GN AVDD 0.072536f
C3 BULKP AVDD 0.120582f
C4 BULKP GNG -0.056171f
C5 BULKP GN -0.16538f
C6 C GN 0.105655f
C7 C BULKP -0.234337f
C8 TIE_H BULKN 0.37082f
C9 MN1/a_324_334# BULKN 0.422f
C10 AVSS BULKN 0.391756f
C11 MN0/a_324_n18# BULKN 0.422415f
C12 AVDD BULKN 0.269584f
C13 GN BULKN 0.410388f
C14 BULKP BULKN 3.595271f
C15 C BULKN 0.568156f
C16 MP1/a_216_334# BULKN 0.091338f
C17 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARBSSW_CV VI CK CKN TIE_L VO1 VO2 XA3/B M4/G AVDD XA4/GNG AVSS
XM1 VI M4/G VO1 AVSS M1/a_324_n18# M2/a_324_n18# SUNSAR_NCHDLR
XM2 VI M4/G VO1 AVSS M2/a_324_n18# M3/a_324_n18# SUNSAR_NCHDLR
XM4 VI M4/G VO1 AVSS M4/a_324_n18# M5/a_324_n18# SUNSAR_NCHDLR
XM3 VI M4/G VO1 AVSS M3/a_324_n18# M4/a_324_n18# SUNSAR_NCHDLR
XM5 VI TIE_L VO2 AVSS M5/a_324_n18# M6/a_324_n18# SUNSAR_NCHDLR
XXCAPB1 XA3/B AVSS XA4/GNG SUNSAR_CAP_BSSW5_CV
XM6 VI TIE_L VO2 AVSS M6/a_324_n18# M7/a_324_n18# SUNSAR_NCHDLR
XM7 VI TIE_L VO2 AVSS M7/a_324_n18# M8/a_324_n18# SUNSAR_NCHDLR
XM8 VI TIE_L VO2 AVSS M8/a_324_n18# M8/a_324_334# SUNSAR_NCHDLR
XXA0 AVDD AVSS CKN AVSS XA0/MP0/a_216_n18# XA3/MP0/a_216_n18# AVDD CK XA0/MN0/a_324_n18#
+ XA3/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA1 XA1/Y AVDD AVDD AVSS AVSS XA4/MP1/a_216_334# XA7/MP1/a_216_n18# XA1/MP0/G XA4/MN1/a_324_334#
+ XA7/MN1/a_324_n18# SUNSAR_TIEH_CV
XXA2 AVDD AVDD AVSS AVSS TIE_L XA7/MP1/a_216_334# XA5/MP1/a_216_n18# XA2/MP0/G XA7/MN1/a_324_334#
+ XA5/MN1/a_324_n18# SUNSAR_TIEL_CV
XXA3 AVDD AVSS AVDD XA4/MN0/a_324_n18# XA3/MP0/S XA3/B XA3/MP0/a_216_n18# VI AVSS
+ CKN XA4/MP0/a_216_n18# XA3/MN0/a_324_n18# SUNSAR_TGPD_CV
XXA5 AVSS XA5/MN1/a_324_n18# XA5/MN1/a_324_334# XA5/MP1/a_216_334# XA5/MP1/a_216_n18#
+ AVDD SUNSAR_TAPCELLB_CV
XXA4 M4/G XA4/GNG XA1/Y AVDD AVSS XA4/MN1/a_324_334# CKN AVDD AVSS XA4/MP0/a_216_n18#
+ XA4/MP1/a_216_334# XA4/MN0/a_324_n18# SUNSAR_SARBSSWCTRL_CV
XXA5b AVSS XA5b/MN1/a_324_n18# XA0/MN0/a_324_n18# XA0/MP0/a_216_n18# XA5b/MP1/a_216_n18#
+ AVDD SUNSAR_TAPCELLB_CV
XXA7 AVSS XA7/MN1/a_324_n18# XA7/MN1/a_324_334# XA7/MP1/a_216_334# XA7/MP1/a_216_n18#
+ AVDD SUNSAR_TAPCELLB_CV
C0 CKN AVDD 0.386132f
C1 AVDD XA0/MP0/a_216_n18# -0.310671f
C2 XA3/MP0/a_216_n18# AVDD -0.316045f
C3 XA7/MP1/a_216_n18# AVDD -0.314169f
C4 M4/G CKN 0.164954f
C5 VI CKN 0.158203f
C6 AVDD XA3/B 1.164377f
C7 XA4/GNG CKN 0.133189f
C8 AVDD XA1/Y 0.335551f
C9 VI XA3/MP0/S 0.083601f
C10 XA4/GNG XA3/B 0.074607f
C11 AVDD XA4/MP0/a_216_n18# -0.315133f
C12 CKN CK 0.081692f
C13 M4/G XA1/Y 0.191529f
C14 XA4/MP1/a_216_334# AVDD -0.311049f
C15 CKN XA3/B 0.220083f
C16 XA1/MP0/G XA1/Y 0.210055f
C17 CKN XA3/MP0/S 0.35416f
C18 XA2/MP0/G AVDD 0.154589f
C19 TIE_L VO2 0.067503f
C20 M4/G VO1 0.121685f
C21 XA4/GNG AVDD 2.419111f
C22 VI VO2 0.402189f
C23 VI VO1 0.51157f
C24 VI TIE_L 0.431984f
C25 VI M4/G 0.734411f
C26 CKN XA1/Y 0.083971f
C27 XA5/MP1/a_216_n18# AVDD -0.312114f
C28 XA7/MP1/a_216_334# AVDD -0.31194f
C29 TIE_L XA2/MP0/G 0.059272f
C30 M4/G XA4/GNG 0.159547f
C31 XA7/MN1/a_324_n18# AVSS 0.352854f
C32 XA5b/MN1/a_324_n18# AVSS 0.422415f
C33 XA0/MN0/a_324_n18# AVSS 0.355076f
C34 AVDD AVSS 16.186546f
C35 XA5b/MP1/a_216_n18# AVSS 0.091271f
C36 XA1/Y AVSS 0.964136f
C37 XA4/MN1/a_324_334# AVSS 0.352614f
C38 XA4/MN0/a_324_n18# AVSS 0.353766f
C39 XA5/MN1/a_324_334# AVSS 0.431299f
C40 XA5/MP1/a_216_334# AVSS 0.091432f
C41 XA3/B AVSS 54.425087f
C42 XA3/MP0/S AVSS 0.743072f
C43 XA7/MN1/a_324_334# AVSS 0.356024f
C44 XA5/MN1/a_324_n18# AVSS 0.354714f
C45 XA2/MP0/G AVSS 0.750734f
C46 XA1/MP0/G AVSS 0.875146f
C47 XA3/MN0/a_324_n18# AVSS 0.351448f
C48 CK AVSS 0.534205f
C49 CKN AVSS 2.229387f
C50 M8/a_324_n18# AVSS 0.354539f
C51 M8/a_324_334# AVSS 0.435553f
C52 M7/a_324_n18# AVSS 0.353892f
C53 VO2 AVSS 0.432698f
C54 TIE_L AVSS 2.998902f
C55 XA4/GNG AVSS 53.063145f
C56 M6/a_324_n18# AVSS 0.353868f
C57 M3/a_324_n18# AVSS 0.353838f
C58 M4/a_324_n18# AVSS 0.353838f
C59 M5/a_324_n18# AVSS 0.355864f
C60 M2/a_324_n18# AVSS 0.353838f
C61 VO1 AVSS 0.482601f
C62 M4/G AVSS 3.126676f
C63 VI AVSS 1.706923f
C64 M1/a_324_n18# AVSS 0.42462f
.ends

.subckt SUNSAR_SAREMX1_CV B EN ENO MP3/a_216_334# MN3/a_324_334# MP3/G A MN2/S BULKP
+ MP0/a_216_n18# AVSS BULKN AVDD RST_N MN0/a_324_n18#
XMP0 AVDD RST_N MP3/G BULKP BULKN MP0/a_216_n18# MP1/a_216_n18# SUNSAR_PCHDL
XMP1 MP2/S B ENO BULKP BULKN MP1/a_216_n18# MP2/a_216_n18# SUNSAR_PCHDL
XMP2 MP3/S A MP2/S BULKP BULKN MP2/a_216_n18# MP3/a_216_n18# SUNSAR_PCHDL
XMN0 MN2/S EN MP3/G BULKN MN0/a_324_n18# MN1/a_324_n18# SUNSAR_NCHDL
XMP3 AVDD MP3/G MP3/S BULKP BULKN MP3/a_216_n18# MP3/a_216_334# SUNSAR_PCHDL
XMN1 MN2/S B AVSS BULKN MN1/a_324_n18# MN2/a_324_n18# SUNSAR_NCHDL
XMN2 AVSS A MN2/S BULKN MN2/a_324_n18# MN3/a_324_n18# SUNSAR_NCHDL
XMN3 ENO MP3/G AVSS BULKN MN3/a_324_n18# MN3/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.236533f
C1 BULKP A 0.108551f
C2 ENO AVSS 0.066248f
C3 MP3/S MP3/G 0.063428f
C4 BULKP B 0.113772f
C5 AVDD AVSS 0.1609f
C6 ENO MP3/G 0.133485f
C7 B A 0.058881f
C8 MP2/S MP3/G 0.064105f
C9 BULKP AVSS 0.059049f
C10 AVDD MP3/G 0.126944f
C11 BULKP MP3/a_216_n18# -0.311038f
C12 RST_N MP3/G 0.054556f
C13 BULKP MP3/G 0.480172f
C14 MP3/G A 0.105132f
C15 ENO MP3/S 0.064105f
C16 MP3/G AVSS 0.051789f
C17 MN2/S AVSS 0.209753f
C18 AVDD MP3/S 0.068807f
C19 MP2/S ENO 0.064105f
C20 BULKP MP2/a_216_n18# -0.311038f
C21 AVDD ENO 0.156546f
C22 AVDD MP2/S 0.055949f
C23 BULKP ENO 0.182005f
C24 BULKP MP1/a_216_n18# -0.311038f
C25 MN3/a_324_n18# BULKN 0.35253f
C26 MN3/a_324_334# BULKN 0.422f
C27 A BULKN 0.498033f
C28 MN2/a_324_n18# BULKN 0.352522f
C29 B BULKN 0.513991f
C30 MN1/a_324_n18# BULKN 0.352522f
C31 AVSS BULKN 0.703356f
C32 MP3/a_216_334# BULKN 0.091338f
C33 MP3/G BULKN 0.827536f
C34 EN BULKN 0.386445f
C35 MN2/S BULKN 0.207484f
C36 MN0/a_324_n18# BULKN 0.422415f
C37 ENO BULKN 0.246284f
C38 AVDD BULKN 0.397419f
C39 BULKP BULKN 7.539519f
C40 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARLTX1_CV RST_N EN LCK_N AVSS MN2/a_324_334# A BULKP MP0/a_216_n18#
+ CHL BULKN AVDD MP2/a_216_334# MN0/a_324_n18#
XMP0 MP1/S RST_N AVDD BULKP BULKN MP0/a_216_n18# RST_N SUNSAR_PCHDL
XMP1 MP2/S RST_N MP1/S BULKP BULKN RST_N RST_N SUNSAR_PCHDL
XMN0 MN1/S A AVSS BULKN MN0/a_324_n18# LCK_N SUNSAR_NCHDL
XMP2 CHL RST_N MP2/S BULKP BULKN RST_N MP2/a_216_334# SUNSAR_PCHDL
XMN1 MN2/S LCK_N MN1/S BULKN A EN SUNSAR_NCHDL
XMN2 CHL EN MN2/S BULKN LCK_N MN2/a_324_334# SUNSAR_NCHDL
C0 AVDD AVSS 0.090662f
C1 AVDD BULKP 0.145188f
C2 MP1/S BULKP -0.050867f
C3 BULKP MP2/S -0.050867f
C4 BULKP RST_N -1.319845f
C5 BULKP CHL 0.074842f
C6 EN BULKN 0.372036f
C7 MN2/a_324_334# BULKN 0.422f
C8 LCK_N BULKN 0.335836f
C9 AVSS BULKN 0.43526f
C10 RST_N BULKN 0.123012f
C11 CHL BULKN 0.260933f
C12 BULKP BULKN 4.387078f
C13 MP2/a_216_334# BULKN 0.091338f
C14 A BULKN 0.372036f
C15 MN0/a_324_n18# BULKN 0.422415f
C16 AVDD BULKN 0.283558f
C17 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARMRYX1_CV CMP_OP CHL_OP CHL_ON XA1/MP3/G RST_N XA5/MP2/a_216_334#
+ ENO XA5/MN2/a_324_334# XA1/MN2/S CMP_ON AVDD AVSS XA2/Y EN
XXA0 AVSS XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ AVDD SUNSAR_TAPCELLB_CV
XXA1 CMP_ON EN ENO XA2/MP0/a_216_n18# XA2/MN0/a_324_n18# XA1/MP3/G CMP_OP XA1/MN2/S
+ AVDD XA1/MP0/a_216_n18# AVSS AVSS AVDD RST_N XA1/MN0/a_324_n18# SUNSAR_SAREMX1_CV
XXA2 AVDD AVSS XA2/Y AVSS XA2/MP0/a_216_n18# XA4/MP0/a_216_n18# AVDD ENO XA2/MN0/a_324_n18#
+ XA4/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA4 RST_N EN XA2/Y AVSS XA5/MN0/a_324_n18# CMP_OP AVDD XA4/MP0/a_216_n18# CHL_OP
+ AVSS AVDD XA5/MP0/a_216_n18# XA4/MN0/a_324_n18# SUNSAR_SARLTX1_CV
XXA5 RST_N EN XA2/Y AVSS XA5/MN2/a_324_334# CMP_ON AVDD XA5/MP0/a_216_n18# CHL_ON
+ AVSS AVDD XA5/MP2/a_216_334# XA5/MN0/a_324_n18# SUNSAR_SARLTX1_CV
C0 AVDD XA2/MP0/a_216_n18# -0.314158f
C1 EN CMP_OP 0.196887f
C2 AVDD XA2/Y 0.086633f
C3 XA2/Y CMP_OP 0.183507f
C4 EN CMP_ON 0.54292f
C5 ENO CMP_OP 0.15365f
C6 XA2/Y CMP_ON 0.130187f
C7 XA2/Y EN 0.114038f
C8 ENO XA1/MP3/G 0.074928f
C9 AVDD RST_N 1.197074f
C10 AVDD CHL_OP 0.06932f
C11 ENO XA2/Y 0.081815f
C12 XA1/MP0/a_216_n18# AVDD -0.312114f
C13 CMP_ON CMP_OP 0.054599f
C14 AVDD XA4/MP0/a_216_n18# -0.314158f
C15 XA1/MP3/G RST_N 0.080501f
C16 AVDD XA5/MP0/a_216_n18# -0.314158f
C17 XA5/MN2/a_324_334# AVSS 0.422f
C18 CHL_ON AVSS 0.232377f
C19 XA5/MP2/a_216_334# AVSS 0.091271f
C20 XA5/MN0/a_324_n18# AVSS 0.353572f
C21 RST_N AVSS 0.223454f
C22 CHL_OP AVSS 0.170116f
C23 XA4/MN0/a_324_n18# AVSS 0.353572f
C24 XA2/MN0/a_324_n18# AVSS 0.353587f
C25 XA2/Y AVSS 1.192111f
C26 XA1/MN3/a_324_n18# AVSS 0.352733f
C27 CMP_OP AVSS 1.304227f
C28 XA1/MN2/a_324_n18# AVSS 0.353381f
C29 CMP_ON AVSS 1.822234f
C30 XA1/MN1/a_324_n18# AVSS 0.358f
C31 XA1/MP3/G AVSS 0.88567f
C32 EN AVSS 2.426762f
C33 XA1/MN2/S AVSS 0.199983f
C34 XA1/MN0/a_324_n18# AVSS 0.35614f
C35 ENO AVSS 0.833836f
C36 XA0/MN1/a_324_n18# AVSS 0.422415f
C37 AVDD AVSS 17.172226f
C38 XA0/MP1/a_216_n18# AVSS 0.091271f
.ends

.subckt SUNSAR_SWX4_CV MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18# Y BULKN
+ AVSS A MN0/a_324_n18# VREF
XMP0 Y A VREF BULKP BULKN MP0/a_216_n18# A SUNSAR_PCHDL
XMP1 VREF A Y BULKP BULKN A A SUNSAR_PCHDL
XMP2 Y A VREF BULKP BULKN A A SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# A SUNSAR_NCHDL
XMP3 VREF A Y BULKP BULKN A MP3/a_216_334# SUNSAR_PCHDL
XMN1 AVSS A Y BULKN A A SUNSAR_NCHDL
XMN2 Y A AVSS BULKN A A SUNSAR_NCHDL
XMN3 AVSS A Y BULKN A MN3/a_324_334# SUNSAR_NCHDL
C0 BULKP VREF 0.287826f
C1 BULKP A -1.606473f
C2 VREF AVSS 0.059626f
C3 A AVSS 0.077171f
C4 Y AVSS 0.183147f
C5 BULKP AVSS 0.063124f
C6 A VREF 0.185495f
C7 Y VREF 0.134317f
C8 Y A 0.147007f
C9 AVSS BULKN 0.671458f
C10 MN3/a_324_334# BULKN 0.422f
C11 MP3/a_216_334# BULKN 0.091338f
C12 VREF BULKN 0.508545f
C13 A BULKN 2.06236f
C14 Y BULKN 0.278638f
C15 MN0/a_324_n18# BULKN 0.422415f
C16 BULKP BULKN 5.176431f
C17 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARCEX1_CV B Y RST AVDD AVSS MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18#
+ BULKN A MN0/a_324_n18#
XMP0 MP1/S A Y BULKP BULKN MP0/a_216_n18# A SUNSAR_PCHDL
XMP1 AVDD A MP1/S BULKP BULKN A B SUNSAR_PCHDL
XMP2 MP3/S B AVDD BULKP BULKN A B SUNSAR_PCHDL
XMN0 MN1/S RST AVSS BULKN MN0/a_324_n18# RST SUNSAR_NCHDL
XMP3 Y B MP3/S BULKP BULKN B MP3/a_216_334# SUNSAR_PCHDL
XMN1 AVSS RST MN1/S BULKN RST RST SUNSAR_NCHDL
XMN2 MN3/S RST AVSS BULKN RST RST SUNSAR_NCHDL
XMN3 Y RST MN3/S BULKN RST MN3/a_324_334# SUNSAR_NCHDL
C0 AVSS Y 0.131513f
C1 BULKP B -1.00547f
C2 BULKP MP3/S -0.050867f
C3 RST Y 0.072094f
C4 BULKP AVDD 0.116689f
C5 BULKP A -1.005062f
C6 BULKP MP1/S -0.050867f
C7 MN1/S AVSS 0.059266f
C8 Y AVDD 0.078529f
C9 BULKP Y 0.191403f
C10 AVSS AVDD 0.10846f
C11 AVDD BULKN 0.253957f
C12 Y BULKN 0.484249f
C13 MN3/a_324_334# BULKN 0.422f
C14 AVSS BULKN 0.502768f
C15 MP3/a_216_334# BULKN 0.091338f
C16 RST BULKN 1.501372f
C17 MN0/a_324_n18# BULKN 0.422415f
C18 B BULKN 0.072331f
C19 A BULKN 0.072331f
C20 BULKP BULKN 5.174408f
C21 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARDIGEX4_CV CMP_OP CMP_ON CP0 CN0 CN1 CEIN XA1/XA2/Y XA9/B DONE XA1/XA1/MP3/G
+ RST_N XA11/A CEO XA4/A CKS XA2/A ENO XA1/XA1/MN2/S CP1 EN VREF XA9/A XA12/A AVSS
+ AVDD
XXA10 AVDD AVSS XA11/A AVSS XA9/MP1/a_216_334# XA11/MP0/a_216_n18# AVDD XA9/Y XA9/MN1/a_324_334#
+ XA11/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA11 AVSS XA12/MN0/a_324_n18# CEIN AVDD AVSS XA11/MP0/a_216_n18# XA12/A XA12/MP0/a_216_n18#
+ AVDD XA11/A XA11/MN0/a_324_n18# SUNSAR_NRX1_CV
XXA12 AVDD AVSS CEO AVSS XA12/MP0/a_216_n18# XA13/MP1/a_216_n18# AVDD XA12/A XA12/MN0/a_324_n18#
+ XA13/MN1/a_324_n18# SUNSAR_IVX1_CV
XXA13 AVSS XA13/MN1/a_324_n18# XA13/MN1/a_324_334# XA13/MP1/a_216_334# XA13/MP1/a_216_n18#
+ AVDD SUNSAR_TAPCELLB_CV
XXA1 CMP_OP XA4/A XA2/A XA1/XA1/MP3/G RST_N XA2/MP0/a_216_n18# ENO XA2/MN0/a_324_n18#
+ XA1/XA1/MN2/S CMP_ON AVDD AVSS XA1/XA2/Y EN SUNSAR_SARMRYX1_CV
XXA2 XA3/MP0/a_216_n18# XA3/MN0/a_324_n18# AVDD XA2/MP0/a_216_n18# CN1 AVSS AVSS XA2/A
+ XA2/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA3 XA4/MP0/a_216_n18# XA4/MN0/a_324_n18# AVDD XA3/MP0/a_216_n18# CP1 AVSS AVSS CN1
+ XA3/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA5 XA6/MP0/a_216_n18# XA6/MN0/a_324_n18# AVDD XA5/MP0/a_216_n18# CN0 AVSS AVSS CP0
+ XA5/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA4 XA5/MP0/a_216_n18# XA5/MN0/a_324_n18# AVDD XA4/MP0/a_216_n18# CP0 AVSS AVSS XA4/A
+ XA4/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA6 CP1 XA9/B CKS AVDD AVSS XA7/MP0/a_216_n18# XA7/MN0/a_324_n18# AVDD XA6/MP0/a_216_n18#
+ AVSS CN0 XA6/MN0/a_324_n18# SUNSAR_SARCEX1_CV
XXA7 AVDD AVSS XA9/A AVSS XA7/MP0/a_216_n18# XA8/MP0/a_216_n18# AVDD ENO XA7/MN0/a_324_n18#
+ XA8/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA8 AVDD AVSS DONE AVSS XA8/MP0/a_216_n18# XA9/MP0/a_216_n18# AVDD XA9/A XA8/MN0/a_324_n18#
+ XA9/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA9 XA9/Y AVDD AVSS XA9/MN1/a_324_334# XA9/B XA9/A AVDD AVSS XA9/MP0/a_216_n18# XA9/MP1/a_216_334#
+ XA9/MN0/a_324_n18# SUNSAR_NDX1_CV
C0 XA2/A CN1 0.328523f
C1 XA9/Y XA9/B 0.108031f
C2 AVDD XA4/A 0.106811f
C3 XA7/MP0/a_216_n18# AVDD -0.312115f
C4 ENO XA9/B 0.051732f
C5 AVDD XA2/MP0/a_216_n18# -0.305873f
C6 AVDD VREF 2.333421f
C7 ENO CMP_ON 0.067952f
C8 XA9/A XA9/B 0.245863f
C9 XA12/A AVDD 0.092808f
C10 ENO CN1 0.083825f
C11 ENO CP1 0.402334f
C12 XA9/Y XA11/A 0.134948f
C13 AVDD XA9/B 0.076896f
C14 AVDD XA5/MP0/a_216_n18# -0.29797f
C15 ENO CP0 0.08098f
C16 XA3/MP0/a_216_n18# AVDD -0.297442f
C17 ENO XA2/A 0.090499f
C18 ENO XA1/XA1/MP3/G 0.086456f
C19 AVDD CN0 0.446492f
C20 VREF XA9/B 0.062419f
C21 CEO AVDD 0.068754f
C22 AVDD CN1 0.116113f
C23 AVDD CP1 0.762798f
C24 CN1 XA4/A 0.465168f
C25 XA12/MP0/a_216_n18# AVDD -0.311437f
C26 CP1 XA4/A 0.193133f
C27 CN0 VREF 0.089615f
C28 AVDD XA8/MP0/a_216_n18# -0.312115f
C29 AVDD CP0 0.188731f
C30 XA11/A AVDD 0.076529f
C31 CP0 XA4/A 0.356664f
C32 AVDD XA2/A 0.204063f
C33 CP1 VREF 1.094435f
C34 XA2/A XA4/A 0.111482f
C35 XA11/MP0/a_216_n18# AVDD -0.31197f
C36 EN XA4/A 0.118846f
C37 XA13/MP1/a_216_n18# AVDD -0.312114f
C38 CEIN XA12/A 0.110841f
C39 XA2/A VREF 0.114185f
C40 CN0 XA9/B 0.069484f
C41 ENO XA9/A 0.07744f
C42 AVDD XA4/MP0/a_216_n18# -0.29797f
C43 XA1/XA2/Y XA4/A 0.161989f
C44 AVDD XA9/MP0/a_216_n18# -0.312114f
C45 XA11/A XA12/A 0.07223f
C46 AVDD XA6/MP0/a_216_n18# -0.305815f
C47 AVDD ENO 2.512355f
C48 ENO XA4/A 0.119363f
C49 CP1 CN0 0.321515f
C50 ENO VREF 0.725442f
C51 DONE XA9/A 0.063409f
C52 CP1 CN1 0.21563f
C53 CP0 CN0 0.301879f
C54 AVDD XA9/A 0.068846f
C55 ENO RST_N 0.661116f
C56 AVDD XA9/MP1/a_216_334# -0.312036f
C57 CP0 CP1 0.177099f
C58 AVDD DONE 0.055251f
C59 XA9/MN1/a_324_334# AVSS 0.355024f
C60 XA9/MN0/a_324_n18# AVSS 0.353772f
C61 XA9/A AVSS 1.385544f
C62 DONE AVSS 0.144723f
C63 XA7/MN0/a_324_n18# AVSS 0.35459f
C64 XA8/MN0/a_324_n18# AVSS 0.355024f
C65 XA9/B AVSS 1.505008f
C66 CKS AVSS 1.45158f
C67 XA6/MN0/a_324_n18# AVSS 0.35614f
C68 XA4/A AVSS 3.135887f
C69 XA4/MN0/a_324_n18# AVSS 0.355615f
C70 CP0 AVSS 2.549277f
C71 CN0 AVSS 0.339688f
C72 XA5/MN0/a_324_n18# AVSS 0.355024f
C73 CN1 AVSS 2.518541f
C74 CP1 AVSS 0.530389f
C75 XA3/MN0/a_324_n18# AVSS 0.355024f
C76 VREF AVSS 0.839587f
C77 XA2/A AVSS 2.066311f
C78 XA2/MN0/a_324_n18# AVSS 0.355615f
C79 XA1/XA5/MN0/a_324_n18# AVSS 0.359841f
C80 RST_N AVSS 0.189551f
C81 XA1/XA4/MN0/a_324_n18# AVSS 0.360407f
C82 XA1/XA2/MN0/a_324_n18# AVSS 0.360407f
C83 XA1/XA2/Y AVSS 1.04564f
C84 XA1/XA1/MN3/a_324_n18# AVSS 0.355196f
C85 CMP_OP AVSS 1.158637f
C86 XA1/XA1/MN2/a_324_n18# AVSS 0.355196f
C87 CMP_ON AVSS 1.344542f
C88 XA1/XA1/MN1/a_324_n18# AVSS 0.355196f
C89 XA1/XA1/MP3/G AVSS 0.827195f
C90 EN AVSS 2.111692f
C91 XA1/XA1/MN2/S AVSS 0.200627f
C92 XA1/XA1/MN0/a_324_n18# AVSS 0.360407f
C93 ENO AVSS 1.876661f
C94 XA1/XA0/MN1/a_324_n18# AVSS 0.422415f
C95 AVDD AVSS 49.990154f
C96 XA1/XA0/MP1/a_216_n18# AVSS 0.091271f
C97 XA13/MN1/a_324_334# AVSS 0.422f
C98 XA13/MP1/a_216_334# AVSS 0.091271f
C99 XA12/MN0/a_324_n18# AVSS 0.355339f
C100 XA13/MN1/a_324_n18# AVSS 0.35614f
C101 CEO AVSS 0.198999f
C102 XA12/A AVSS 0.873459f
C103 XA11/MN0/a_324_n18# AVSS 0.355024f
C104 CEIN AVSS 0.470328f
C105 XA11/A AVSS 0.773929f
C106 XA9/Y AVSS 0.833236f
.ends

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW
+ VREF AVDD AVSS
*.subckt SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4> D<3>
*+ D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
XXDAC1 XA0/CP0 D<7> XA1/CP0 D<6> XA2/CP0 D<5> XA3/CP0 D<4> D<3> D<2> D<1> SARP XDAC1/XC1/XRES1A/B
+ XA0/CP1 AVSS AVSS SUNSAR_CDAC8_CV
XXDAC2 XA0/CN0 XA1/CN1 XA1/CN0 XA2/CN1 XA2/CN0 XA3/CN1 XA3/CN0 XA4/CN0 XA5/CN0 XA6/CN0
+ XA7/CN0 SARN XDAC2/XC1/XRES1A/B D<8> AVSS AVSS SUNSAR_CDAC8_CV
XXA20 SARP SARN XA8/CEO XA20/XA12/Y XA20/XA3/CO XA20/XA3a/A CK_SAMPLE XA20/XA9/A XA20/CPO
+ DONE AVSS XA20/CNO AVDD SUNSAR_SARCMPX1_CV
XXB1 SAR_IP CK_SAMPLE_BSSW XB1/CKN XA0/CEIN SARP SARN XB1/XA3/B XB1/M4/G AVDD XB1/XA4/GNG
+ AVSS SUNSAR_SARBSSW_CV
XXA0 XA20/CPO XA20/CNO XA0/CP0 XA0/CN0 D<8> XA0/CEIN XA0/XA1/XA2/Y XA0/XA9/B XA0/DONE
+ XA0/XA1/XA1/MP3/G EN XA0/XA11/A XA0/CEO XA0/XA4/A CK_SAMPLE XA0/XA2/A XA1/EN XA0/XA1/XA1/MN2/S
+ XA0/CP1 EN VREF XA0/XA9/A XA0/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA1 XA20/CPO XA20/CNO XA1/CP0 XA1/CN0 XA1/CN1 XA0/CEO XA1/XA1/XA2/Y XA1/XA9/B XA1/DONE
+ XA1/XA1/XA1/MP3/G EN XA1/XA11/A XA1/CEO XA1/XA4/A CK_SAMPLE XA1/XA2/A XA2/EN XA1/XA1/XA1/MN2/S
+ D<7> XA1/EN VREF XA1/XA9/A XA1/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXB2 SAR_IN CK_SAMPLE_BSSW XB2/CKN XA0/CEIN SARN SARP XB2/XA3/B XB2/M4/G AVDD XB2/XA4/GNG
+ AVSS SUNSAR_SARBSSW_CV
XXA2 XA20/CPO XA20/CNO XA2/CP0 XA2/CN0 XA2/CN1 XA1/CEO XA2/XA1/XA2/Y XA2/XA9/B XA2/DONE
+ XA2/XA1/XA1/MP3/G EN XA2/XA11/A XA2/CEO XA2/XA4/A CK_SAMPLE XA2/XA2/A XA3/EN XA2/XA1/XA1/MN2/S
+ D<6> XA2/EN VREF XA2/XA9/A XA2/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA3 XA20/CPO XA20/CNO XA3/CP0 XA3/CN0 XA3/CN1 XA2/CEO XA3/XA1/XA2/Y XA3/XA9/B XA3/DONE
+ XA3/XA1/XA1/MP3/G EN XA3/XA11/A XA3/CEO XA3/XA4/A CK_SAMPLE XA3/XA2/A XA4/EN XA3/XA1/XA1/MN2/S
+ D<5> XA3/EN VREF XA3/XA9/A XA3/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA4 XA20/CPO XA20/CNO XA4/CP0 XA4/CN0 XA4/CN1 XA3/CEO XA4/XA1/XA2/Y XA4/XA9/B XA4/DONE
+ XA4/XA1/XA1/MP3/G EN XA4/XA11/A XA4/CEO XA4/XA4/A CK_SAMPLE XA4/XA2/A XA5/EN XA4/XA1/XA1/MN2/S
+ D<4> XA4/EN VREF XA4/XA9/A XA4/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA5 XA20/CPO XA20/CNO XA5/CP0 XA5/CN0 XA5/CN1 XA4/CEO XA5/XA1/XA2/Y XA5/XA9/B XA5/DONE
+ XA5/XA1/XA1/MP3/G EN XA5/XA11/A XA5/CEO XA5/XA4/A CK_SAMPLE XA5/XA2/A XA6/EN XA5/XA1/XA1/MN2/S
+ D<3> XA5/EN VREF XA5/XA9/A XA5/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA6 XA20/CPO XA20/CNO XA6/CP0 XA6/CN0 XA6/CN1 XA5/CEO XA6/XA1/XA2/Y XA6/XA9/B XA6/DONE
+ XA6/XA1/XA1/MP3/G EN XA6/XA11/A XA6/CEO XA6/XA4/A CK_SAMPLE XA6/XA2/A XA7/EN XA6/XA1/XA1/MN2/S
+ D<2> XA6/EN VREF XA6/XA9/A XA6/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA7 XA20/CPO XA20/CNO XA7/CP0 XA7/CN0 XA7/CN1 XA6/CEO XA7/XA1/XA2/Y XA7/XA9/B XA7/DONE
+ XA7/XA1/XA1/MP3/G EN XA7/XA11/A XA7/CEO XA7/XA4/A CK_SAMPLE XA7/XA2/A XA8/EN XA7/XA1/XA1/MN2/S
+ D<1> XA7/EN VREF XA7/XA9/A XA7/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA8 XA20/CPO XA20/CNO XA8/CP0 XA8/CN0 XA8/CN1 XA7/CEO XA8/XA1/XA2/Y XA8/XA9/B DONE
+ XA8/XA1/XA1/MP3/G EN XA8/XA11/A XA8/CEO XA8/XA4/A CK_SAMPLE XA8/XA2/A XA8/ENO XA8/XA1/XA1/MN2/S
+ D<0> XA8/EN VREF XA8/XA9/A XA8/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
C0 XA20/CNO XA8/XA4/A 0.141687f
C1 XA1/CN1 XA0/CN0 0.588325f
C2 EN XA6/XA4/A 0.088464f
C3 EN XA1/CN1 0.097358f
C4 CK_SAMPLE XA8/EN 0.09249f
C5 XA3/CN1 XA0/CN0 0.068528f
C6 XA3/CN0 D<3> 0.128372f
C7 EN XA3/CN1 0.09808f
C8 CK_SAMPLE XA5/XA9/B 0.078536f
C9 XA5/XA4/A XA6/XA4/A 0.082663f
C10 AVDD XA4/EN 0.091274f
C11 D<5> XA0/CN0 0.055822f
C12 XA4/CEO XA5/XA12/A 0.084465f
C13 EN D<5> 0.064647f
C14 XA1/CN1 XA0/CP1 1.772852f
C15 XA1/EN XA20/CPO 0.251162f
C16 VREF XA0/CN0 0.072034f
C17 XA20/CNO D<6> 0.055536f
C18 XA20/CPO XA4/XA1/XA2/Y 0.069955f
C19 XA2/CN1 D<4> 0.066149f
C20 XA1/CEO XA1/XA12/A 0.264747f
C21 EN VREF 0.820466f
C22 XA7/CN0 XA6/CN0 2.515831f
C23 D<7> D<8> 0.073351f
C24 CK_SAMPLE D<2> 0.100705f
C25 XA3/CN1 XA0/CP1 0.145077f
C26 EN XA7/EN 0.311924f
C27 XA2/EN EN 0.235384f
C28 XA1/CP0 XA2/CN1 0.138993f
C29 XA1/CN1 XA4/CN0 0.072536f
C30 XA5/CN0 XA6/CN0 1.602954f
C31 XB1/XA4/GNG SARP 1.731831f
C32 D<1> D<8> 0.077821f
C33 XA0/XA4/A EN 0.080713f
C34 D<2> XA1/CN0 0.079442f
C35 D<5> XA0/CP1 0.397308f
C36 XA2/CN1 XA1/CN0 0.547568f
C37 AVDD XA3/EN 0.792171f
C38 SARN XB1/M4/G 0.156054f
C39 XA2/CEO AVDD 1.281467f
C40 XA0/CP0 XA0/CN0 5.679079f
C41 XA3/CN1 XA4/CN0 0.066873f
C42 AVDD XA4/CP0 -0.059324f
C43 EN XA0/CP0 0.063812f
C44 D<4> D<3> 0.673295f
C45 VREF XA0/CP1 0.083267f
C46 XA20/CNO XA6/CN0 0.062575f
C47 AVDD XA3/CEO 0.346649f
C48 XA8/XA9/A DONE 0.099743f
C49 XA2/CN0 XA6/CN0 0.090965f
C50 CK_SAMPLE D<3> 0.1008f
C51 XA20/CNO XA2/CP0 0.057246f
C52 XA2/CN0 XA2/CP0 2.959908f
C53 XA1/XA4/A XA2/XA4/A 0.082663f
C54 VREF XA4/CN0 0.072034f
C55 D<3> XA1/CN0 0.095342f
C56 VREF XA5/EN 0.153675f
C57 XA3/EN XA4/EN 1.263078f
C58 EN XA8/XA2/A 0.11426f
C59 SARN XA20/XA9/A 0.426703f
C60 XA2/CP0 XA3/CP0 0.876237f
C61 XA20/CPO XA1/CN1 0.26688f
C62 XA0/CP0 XA0/CP1 3.663675f
C63 XA3/CN0 XA6/CN0 0.066517f
C64 CK_SAMPLE XA4/XA9/B 0.07743f
C65 SAR_IP XA0/CEIN 0.064942f
C66 XA20/CPO XA3/CN1 0.273087f
C67 AVDD XA0/CN0 3.027888f
C68 XB2/XA4/GNG XDAC2/XC1/XRES16/B 0.098205f
C69 AVDD EN 3.259237f
C70 EN XA7/XA4/A 0.088236f
C71 XA2/CN1 D<2> 0.065888f
C72 XA20/CPO D<5> 0.063761f
C73 CK_SAMPLE D<6> 0.100705f
C74 XA1/EN XA20/CNO 0.302764f
C75 XA0/CN0 D<8> 0.492996f
C76 AVDD SARN 0.121416f
C77 EN D<8> 0.331359f
C78 XA1/CP0 D<6> 0.994598f
C79 XA5/XA11/A XA4/CEO 0.06726f
C80 XA20/CNO XA2/XA4/A 0.212165f
C81 D<6> XA1/CN0 0.063251f
C82 XA2/CEO XA3/CEO 0.431792f
C83 XA1/XA4/A XA1/CN1 0.092714f
C84 XA20/CPO XA7/EN 0.251162f
C85 XA2/EN XA20/CPO 0.378571f
C86 SARN D<8> 0.061494f
C87 D<7> XA0/CN0 0.055917f
C88 EN XA4/EN 0.235384f
C89 D<3> D<2> 1.425882f
C90 XA2/CN1 D<3> 0.066027f
C91 EN D<7> 0.064647f
C92 XA3/CN1 SARP 0.06043f
C93 VREF XA6/EN 0.153675f
C94 CK_SAMPLE XA6/CN0 0.070742f
C95 XA1/CN1 XA7/CN0 0.076884f
C96 XA20/CPO XA0/CP0 0.060601f
C97 XA2/CP0 D<4> 0.22346f
C98 D<1> XA0/CN0 0.182038f
C99 XA0/CP1 D<8> 0.794747f
C100 EN XA6/XA2/A 0.11426f
C101 AVDD XA4/CN0 3.073464f
C102 EN D<1> 0.072042f
C103 AVDD XA5/EN 0.79217f
C104 XA3/CN1 XA7/CN0 0.070443f
C105 XB2/M4/G XA0/CEIN 0.131052f
C106 XA1/CN1 XA5/CN0 0.072507f
C107 XA1/XA2/A EN 0.11418f
C108 XA6/CN0 XA1/CN0 0.086627f
C109 XA1/CP0 XA2/CP0 0.543831f
C110 D<7> XA0/CP1 0.09073f
C111 XA4/CN0 D<8> 0.073409f
C112 XA2/CP0 XA1/CN0 0.064892f
C113 EN XA3/EN 0.311923f
C114 XB1/M4/G SARP 0.145435f
C115 XA20/CNO XA6/XA4/A 0.212165f
C116 XA3/CN1 XA5/CN0 0.066278f
C117 XA20/CNO XA1/CN1 0.19049f
C118 XA1/CN1 XA2/CN0 0.079559f
C119 XB1/XA4/GNG XDAC1/XC1/XRES1A/B 0.403704f
C120 VREF XA7/CN0 0.074599f
C121 D<6> XA2/CN1 0.418934f
C122 AVDD CK_SAMPLE_BSSW 18.810143f
C123 XA20/CNO XA3/CN1 0.193771f
C124 XA7/EN XA7/CN0 0.141771f
C125 XA1/CN1 XA3/CP0 0.071833f
C126 XB2/XA4/GNG XDAC2/XC1/XRES1A/B 0.403704f
C127 XA2/CN0 XA3/CN1 0.493041f
C128 XA0/CP0 SARP 0.103942f
C129 SAR_IN SARN 0.279434f
C130 VREF XA5/CN0 0.074599f
C131 AVDD XA20/CPO 3.731571f
C132 XA4/CN0 D<1> 0.073242f
C133 XA5/CN0 XA5/CP0 0.119737f
C134 XA20/CNO D<5> 0.056276f
C135 XA7/CEO XA7/XA11/A 0.126482f
C136 XA1/EN CK_SAMPLE 0.092446f
C137 XA2/CN0 D<5> 0.055822f
C138 XA1/CN1 XA3/CN0 0.075909f
C139 XA3/CN1 XA3/CP0 0.174111f
C140 XA6/CN0 XA6/CN1 0.050253f
C141 CK_SAMPLE DONE 0.117757f
C142 XA20/CPO D<8> 0.223309f
C143 XA1/EN XA1/CP0 0.061526f
C144 XA20/CNO VREF 0.116975f
C145 VREF XA2/CN0 0.072034f
C146 XA3/CN1 XA3/CN0 0.600488f
C147 D<5> XA3/CP0 3.918876f
C148 XA1/EN XA1/CN0 0.058697f
C149 XA6/CN0 D<2> 1.503286f
C150 XA2/CN1 XA6/CN0 0.065942f
C151 XA20/CNO XA7/EN 0.30307f
C152 AVDD XA6/EN 0.091274f
C153 XA5/EN XA5/XA1/XA1/MP3/G 0.095485f
C154 EN XA7/XA2/A 0.11418f
C155 XA2/EN XA20/CNO 0.457819f
C156 EN XA0/CN0 0.067256f
C157 XA20/CPO XA6/XA1/XA2/Y 0.069955f
C158 XA4/CP0 XA4/CN0 0.123858f
C159 AVDD XA5/CEO 0.346649f
C160 XA20/CPO XA4/EN 0.378571f
C161 XA2/CN1 XA2/CP0 0.105717f
C162 XA20/CPO D<7> 0.063761f
C163 D<5> XA3/CN0 0.09973f
C164 XA0/XA4/A XA20/CNO 0.212165f
C165 SARN XA0/CN0 0.105779f
C166 XA2/XA1/XA1/MP3/G XA3/EN 0.058161f
C167 CK_SAMPLE XA3/XA9/B 0.078536f
C168 VREF XA3/CN0 0.074599f
C169 XA20/CNO XA0/CP0 0.057246f
C170 XA6/CEO XA7/CEO 0.431793f
C171 AVDD SARP 0.084261f
C172 XB1/XA4/GNG XDAC1/XC1/XRES16/B 0.098205f
C173 XA20/CPO D<1> 0.072437f
C174 EN XA5/XA4/A 0.088236f
C175 D<3> XA6/CN0 0.152644f
C176 XA6/CP0 XA6/CN0 0.123858f
C177 VREF XA8/ENO 0.141848f
C178 EN XA0/CP1 0.068664f
C179 SARP D<8> 0.204103f
C180 XA3/CP0 XA0/CP0 0.133088f
C181 AVDD XA7/CN0 3.327564f
C182 XA1/CN1 D<4> 0.107054f
C183 XA20/CPO XA3/EN 0.251162f
C184 XA4/CN0 XA0/CN0 0.073539f
C185 XA3/CN1 D<4> 0.249488f
C186 AVDD XA5/CN0 3.17708f
C187 XA6/CEO XA7/XA12/A 0.084465f
C188 XA7/CN0 D<8> 0.077804f
C189 XA1/CN1 XA1/CP0 0.183042f
C190 EN XA2/XA2/A 0.11426f
C191 EN XA4/CN0 0.071817f
C192 XA1/EN XA0/XA1/XA1/MP3/G 0.058161f
C193 EN XA5/EN 0.311924f
C194 XA20/CNO XA20/XA3a/A 0.092122f
C195 XA1/CN1 XA1/CN0 0.71203f
C196 D<5> D<4> 0.103559f
C197 XA1/CP0 XA3/CN1 0.13878f
C198 XA2/CN1 XA2/XA4/A 0.064665f
C199 XA5/CN0 D<8> 0.073351f
C200 VREF XA6/CEO 0.367402f
C201 AVDD XA20/CNO 3.58161f
C202 XA20/CNO XA7/XA4/A 0.286188f
C203 CK_SAMPLE D<5> 0.1008f
C204 AVDD XA2/CN0 3.034707f
C205 XA3/CN1 XA1/CN0 0.068986f
C206 VREF D<4> 0.083267f
C207 XA1/CP0 D<5> 0.133712f
C208 CK_SAMPLE VREF 2.128126f
C209 XA20/CNO D<8> 0.179623f
C210 D<5> XA1/CN0 0.055822f
C211 AVDD XA3/CP0 0.065787f
C212 D<1> XA7/CN0 2.80043f
C213 XA2/CN0 D<8> 0.078197f
C214 CK_SAMPLE XA7/EN 0.092446f
C215 D<6> XA2/CP0 4.248191f
C216 XA6/EN XA5/XA1/XA1/MN2/S 0.064012f
C217 XA2/EN CK_SAMPLE 0.09249f
C218 XA20/CPO XA0/CN0 0.057021f
C219 VREF XA1/CN0 0.074599f
C220 XA2/CEO XA3/XA12/A 0.084465f
C221 AVDD XA3/CN0 3.158329f
C222 SAR_IN SARP 0.093333f
C223 XA2/EN XA1/CP0 0.092109f
C224 XA20/CPO EN 0.811076f
C225 XA20/CNO XA4/EN 0.457818f
C226 XA3/CP0 D<8> 0.073351f
C227 XA5/CN0 D<1> 0.073281f
C228 XA20/CNO D<7> 0.056276f
C229 XB2/CKN XA0/CEIN 0.064949f
C230 XA3/XA12/A XA3/CEO 0.264747f
C231 XA2/EN XA1/CN0 0.121195f
C232 XA5/EN XA4/CN0 0.060344f
C233 XA3/CN0 D<8> 0.073427f
C234 AVDD XA8/ENO 0.380956f
C235 EN XA4/XA4/A 0.088464f
C236 VREF XA8/EN 0.153676f
C237 XA4/EN XA3/CP0 0.092109f
C238 XA1/CP0 XA0/CP0 2.100499f
C239 XA20/CNO D<1> 0.064523f
C240 XA1/CN1 D<2> 0.104749f
C241 XA1/CN1 XA2/CN1 3.366419f
C242 XA2/CN0 D<1> 0.079819f
C243 EN XA6/EN 0.235384f
C244 XA7/EN XA8/EN 1.263078f
C245 AVDD XB2/XA3/B 0.138847f
C246 XA3/XA4/A XA3/CN1 0.092714f
C247 XA4/EN XA3/CN0 0.121195f
C248 XA20/CPO XA0/CP1 0.062543f
C249 EN XA4/XA2/A 0.11426f
C250 XA3/CN1 D<2> 0.065873f
C251 XA2/CN1 XA3/CN1 1.324099f
C252 XA20/CNO XA3/EN 0.302924f
C253 AVDD XA7/CP0 -0.059568f
C254 XA2/CN0 XA3/EN 0.056267f
C255 CK_SAMPLE D<0> 0.081532f
C256 EN XA1/XA4/A 0.088236f
C257 XA2/CN1 D<5> 0.066437f
C258 AVDD XA6/CEO 1.281468f
C259 XA3/CN0 D<1> 0.076653f
C260 XA20/CPO XA4/CN0 0.064431f
C261 XA20/CPO XA5/XA1/XA2/Y 0.078271f
C262 XA20/CPO XA5/EN 0.251162f
C263 XA1/CN1 D<3> 0.221986f
C264 XA3/EN XA3/CP0 0.061526f
C265 VREF XA0/CEIN 0.057694f
C266 XA2/XA1/XA2/Y XA20/CPO 0.069955f
C267 XA0/CEO XA1/XA11/A 0.06726f
C268 XA20/CPO XA1/XA1/XA2/Y 0.078271f
C269 VREF D<2> 0.083267f
C270 AVDD CK_SAMPLE 4.54462f
C271 XA7/CN0 XA0/CN0 0.078508f
C272 XA0/CEIN XB1/M4/G 0.129829f
C273 SARN SARP 5.580191f
C274 EN XA7/CN0 0.07142f
C275 XA3/EN XA3/CN0 0.058697f
C276 XA3/CN1 D<3> 0.065888f
C277 AVDD XA1/CP0 0.065787f
C278 XA2/EN XA2/CN1 0.336727f
C279 D<4> D<8> 0.073479f
C280 XA5/CN0 XA0/CN0 0.073399f
C281 AVDD XA1/CN0 3.153384f
C282 CK_SAMPLE XA2/XA9/B 0.07743f
C283 XA5/EN XA6/EN 1.263079f
C284 EN XA5/CN0 0.071169f
C285 XA1/CP0 D<8> 0.073351f
C286 XA2/CN1 XA0/CP0 0.133733f
C287 VREF D<3> 0.08346f
C288 XA1/CN0 D<8> 0.079787f
C289 XA20/CNO XA0/CN0 0.055193f
C290 CK_SAMPLE XA4/EN 0.09249f
C291 CK_SAMPLE D<7> 0.1008f
C292 XA20/CNO EN 2.6376f
C293 XA2/CN0 XA0/CN0 0.081585f
C294 AVDD XA8/EN 0.092467f
C295 CK_SAMPLE XA8/XA9/B 0.180961f
C296 EN XA2/CN0 0.065579f
C297 XA1/CP0 D<7> 4.346893f
C298 XA1/CN1 D<6> 0.071041f
C299 XA3/CP0 XA0/CN0 0.127416f
C300 D<7> XA1/CN0 0.099794f
C301 CK_SAMPLE D<1> 0.1008f
C302 VREF XA4/CEO 0.367402f
C303 EN XA3/CP0 0.061409f
C304 XA4/CN0 XA7/CN0 0.097179f
C305 XA20/CNO XA5/XA4/A 0.286129f
C306 D<6> XA3/CN1 0.142972f
C307 XA5/EN XA7/CN0 0.068436f
C308 XA3/CN0 XA0/CN0 0.077181f
C309 XA20/CPO XA6/EN 0.378571f
C310 XA20/CPO XA8/XA1/XA2/Y 0.081818f
C311 EN XA3/CN0 0.064814f
C312 D<1> XA1/CN0 0.07983f
C313 XA20/CNO XA0/CP1 0.055536f
C314 CK_SAMPLE XA3/EN 0.092446f
C315 XA4/CN0 XA5/CN0 1.498409f
C316 D<6> D<5> 0.269031f
C317 XA5/EN XA5/CN0 0.064699f
C318 AVDD XA0/CEIN 12.483942f
C319 XA1/CN1 XA6/CN0 0.072489f
C320 VREF D<6> 0.083267f
C321 CK_SAMPLE XA1/XA9/B 0.078536f
C322 XA20/CNO XA4/CN0 0.062602f
C323 CK_SAMPLE XA6/XA9/B 0.07743f
C324 XA6/XA1/XA1/MP3/G XA7/EN 0.058161f
C325 D<1> XA8/EN 0.096733f
C326 XA1/CN1 XA2/CP0 0.070579f
C327 XA20/CNO XA5/EN 0.302925f
C328 XA2/CN0 XA4/CN0 0.067819f
C329 D<2> D<8> 0.086175f
C330 XA2/CN1 D<8> 0.706063f
C331 XA3/CN1 XA6/CN0 0.066079f
C332 XA7/XA1/XA1/MN2/S XA8/EN 0.064012f
C333 XA20/CPO XA7/CN0 0.063388f
C334 XA2/CP0 XA3/CN1 0.135532f
C335 AVDD XA6/CP0 -0.059324f
C336 D<6> XA0/CP0 0.134985f
C337 XA2/CN1 D<7> 0.14594f
C338 XA2/CP0 D<5> 0.755024f
C339 XA3/CN0 XA4/CN0 1.953506f
C340 XA20/CPO XA5/CN0 0.063388f
C341 VREF XA6/CN0 0.072034f
C342 D<4> XA0/CN0 0.075722f
C343 XA7/XA4/A XA8/XA4/A 0.082663f
C344 EN D<4> 0.071321f
C345 XA20/CPO XA20/XA3/CO 0.314324f
C346 CK_SAMPLE XA0/CN0 0.070742f
C347 XA7/EN XA6/CN0 0.060348f
C348 D<3> D<8> 0.073443f
C349 XB2/XA4/GNG SARN 1.731831f
C350 D<1> D<2> 2.044239f
C351 XA2/CN1 D<1> 0.070327f
C352 XA1/CEO XA1/XA11/A 0.126482f
C353 AVDD XA4/CEO 1.281468f
C354 XA20/CNO XA20/CPO 7.4485f
C355 XA1/CP0 XA0/CN0 0.112242f
C356 XA20/CPO XA2/CN0 0.057021f
C357 EN XA1/CP0 0.061409f
C358 XA1/CN0 XA0/CN0 3.463352f
C359 XA1/EN XA1/CN1 0.231584f
C360 XA5/CN0 XA6/EN 0.13162f
C361 XA2/EN XA1/XA1/XA1/MN2/S 0.064012f
C362 EN XA1/CN0 0.064814f
C363 XA20/CPO XA3/CP0 0.060463f
C364 XA20/CNO XA4/XA4/A 0.212165f
C365 SAR_IN XA0/CEIN 0.069519f
C366 XA2/CP0 XA0/CP0 0.132811f
C367 XA20/CNO XA6/EN 0.457818f
C368 CK_SAMPLE XA0/CP1 0.100695f
C369 XA4/CN1 XA4/CN0 0.050253f
C370 D<1> D<3> 0.155191f
C371 XA20/CPO XA3/CN0 0.055878f
C372 EN XA8/EN 0.235644f
C373 D<4> XA4/CN0 1.354956f
C374 XA1/EN VREF 0.153675f
C375 XA20/CNO XA1/XA4/A 0.286128f
C376 D<6> D<8> 0.073351f
C377 XA20/CPO XA8/ENO 0.12399f
C378 CK_SAMPLE XA4/CN0 0.070742f
C379 XA5/CN0 XA7/CN0 0.076127f
C380 CK_SAMPLE XA5/EN 0.092446f
C381 VREF DONE 0.089716f
C382 XA5/XA12/A XA5/CEO 0.264747f
C383 XA2/EN XA1/EN 1.263076f
C384 XA0/XA2/A EN 0.11426f
C385 XA4/CN0 XA1/CN0 0.06659f
C386 D<6> D<7> 1.431497f
C387 AVDD XA6/CN0 3.046785f
C388 XA20/CNO XA7/CN0 0.061266f
C389 D<2> XA0/CN0 0.092459f
C390 XA2/CN1 XA0/CN0 0.068595f
C391 EN XA3/XA4/A 0.088236f
C392 XA2/CN0 XA7/CN0 0.071338f
C393 EN D<2> 0.071321f
C394 AVDD XA2/CP0 0.056743f
C395 EN XA2/CN1 0.099922f
C396 XA0/CEO VREF 0.367402f
C397 XA20/CNO XA5/CN0 0.060347f
C398 XA7/CEO XA7/XA12/A 0.264746f
C399 XA6/CN0 D<8> 0.073351f
C400 SAR_IP SARN 0.203788f
C401 XA2/CN0 XA5/CN0 0.068349f
C402 SARN XA0/CEIN 0.28158f
C403 XA1/CN1 XA3/CN1 0.071724f
C404 XA20/CPO D<4> 0.071274f
C405 XA20/CNO XA20/XA3/CO 0.129958f
C406 XA2/CP0 D<8> 0.073351f
C407 EN XA3/XA2/A 0.11418f
C408 XA20/CPO XA3/XA1/XA2/Y 0.078271f
C409 XA3/CN0 XA7/CN0 0.071524f
C410 XA1/CN1 D<5> 0.228006f
C411 XA20/CPO XA1/CP0 0.060463f
C412 XA20/CNO XA2/CN0 0.055193f
C413 D<3> XA0/CN0 0.087399f
C414 XA2/CN1 XA0/CP1 0.147379f
C415 EN D<3> 0.072042f
C416 XA2/CP0 D<7> 1.259954f
C417 XA20/CPO XA1/CN0 0.055878f
C418 XA3/CN0 XA5/CN0 0.10727f
C419 D<5> XA3/CN1 0.674953f
C420 CK_SAMPLE XA0/XA9/B 0.07743f
C421 XA20/CNO XA3/CP0 0.056087f
C422 CK_SAMPLE XA7/XA9/B 0.078889f
C423 EN XA8/XA4/A 0.084632f
C424 D<1> XA6/CN0 0.073349f
C425 AVDD XB1/XA3/B 0.138847f
C426 XA2/CN0 XA3/CP0 0.058117f
C427 CK_SAMPLE XA6/EN 0.09249f
C428 VREF XA8/CEO 0.179573f
C429 XA2/EN XA1/CN1 0.109215f
C430 XA4/CN0 D<2> 0.066013f
C431 XA2/CN1 XA4/CN0 0.066079f
C432 AVDD XA1/EN 0.7922f
C433 XA20/CNO XA3/CN0 0.053255f
C434 XA2/CN0 XA3/CN0 1.917195f
C435 XA20/CPO XA8/EN 0.376936f
C436 AVDD DONE 0.873653f
C437 XA8/ENO XA20/XA3/CO 0.159182f
C438 VREF D<5> 0.08346f
C439 XA7/CN0 XA7/CP0 0.119737f
C440 XA1/CN1 XA0/CP0 0.137819f
C441 XA1/CEO XA0/CEO 0.431792f
C442 XA20/CNO XA8/ENO 0.133232f
C443 XA3/CN0 XA3/CP0 2.962606f
C444 XB2/M4/G SARN 0.248185f
C445 XA3/CN1 XA0/CP0 0.147255f
C446 D<6> XA0/CN0 0.056493f
C447 VREF XA7/EN 0.153675f
C448 XA4/CN0 D<3> 0.097821f
C449 CK_SAMPLE XA20/XA12/Y 0.070809f
C450 AVDD XA0/CEO 1.281467f
C451 XA2/EN VREF 0.153675f
C452 EN D<6> 0.063885f
C453 CK_SAMPLE_BSSW XA0/CEIN 7.032176f
C454 CK_SAMPLE XA7/CN0 0.071155f
C455 XA1/EN D<7> 0.063821f
C456 XA5/EN D<3> 0.070845f
C457 XA5/EN XA4/XA1/XA1/MP3/G 0.058161f
C458 D<5> XA0/CP0 0.140102f
C459 XA5/XA11/A XA5/CEO 0.126483f
C460 XA20/CPO D<2> 0.071274f
C461 XA20/CPO XA2/CN1 0.240418f
C462 XB1/CKN XA0/CEIN 0.064949f
C463 CK_SAMPLE XA5/CN0 0.071155f
C464 XA7/CN0 XA1/CN0 0.071267f
C465 AVDD XA7/CEO 0.348648f
C466 XA20/CPO XA7/XA1/XA2/Y 0.078271f
C467 XA20/CNO D<4> 0.064267f
C468 XA3/XA4/A XA4/XA4/A 0.082663f
C469 XA2/CN0 D<4> 0.070487f
C470 XA5/CN0 XA1/CN0 0.066254f
C471 D<6> XA0/CP1 0.129555f
C472 XA6/CN0 XA0/CN0 0.090338f
C473 EN XA6/CN0 0.071885f
C474 CK_SAMPLE XA2/CN0 0.070742f
C475 XA7/CN0 XA8/EN 0.131865f
C476 XA20/CNO XA1/CP0 0.056087f
C477 XA2/CP0 XA0/CN0 0.058178f
C478 XA4/EN XA3/XA1/XA1/MN2/S 0.064012f
C479 AVDD XA8/CEO 1.016913f
C480 XA3/CP0 D<4> 0.861557f
C481 EN XA2/CP0 0.06151f
C482 XA20/CPO D<3> 0.072437f
C483 XA20/CNO XA1/CN0 0.053255f
C484 XA1/CN1 D<8> 0.205177f
C485 VREF D<0> 0.076849f
C486 XA1/XA1/XA1/MP3/G XA1/EN 0.095485f
C487 XA2/CN0 XA1/CN0 2.589554f
C488 SAR_IP SARP 0.285355f
C489 XA3/EN XA3/XA1/XA1/MP3/G 0.095485f
C490 XA3/CN0 D<4> 0.077262f
C491 XA6/CEO XA7/XA11/A 0.06726f
C492 XA1/CP0 XA3/CP0 0.722823f
C493 XA0/CEIN SARP 0.45294f
C494 XA2/CN1 SARP 0.050102f
C495 XA3/CN1 D<8> 1.32017f
C496 CK_SAMPLE XA3/CN0 0.071155f
C497 XA0/CEO XA1/XA12/A 0.084465f
C498 XA3/CP0 XA1/CN0 0.058178f
C499 XA1/CN1 D<7> 0.547462f
C500 AVDD VREF 19.060085f
C501 XA20/CNO XA8/EN 0.455652f
C502 XA6/EN D<3> 0.096733f
C503 D<5> D<8> 0.073541f
C504 AVDD XA5/CP0 -0.059568f
C505 XA3/CN0 XA1/CN0 0.070946f
C506 AVDD XA7/EN 0.792171f
C507 XA7/CN0 D<2> 0.142721f
C508 XA2/CN1 XA7/CN0 0.070367f
C509 CK_SAMPLE XA8/ENO 0.111631f
C510 XA4/EN XA3/CN1 0.112126f
C511 XA2/EN AVDD 0.091274f
C512 XA3/CN1 D<7> 0.139054f
C513 XA1/CN1 D<1> 0.076935f
C514 XA4/CN0 XA6/CN0 0.099672f
C515 XA4/EN D<5> 0.084621f
C516 D<5> D<7> 0.146139f
C517 XA1/EN XA0/CN0 0.056267f
C518 XA5/CN0 D<2> 0.066074f
C519 XA2/CN1 XA5/CN0 0.06599f
C520 XA1/EN EN 0.315014f
C521 XA3/CN1 D<1> 0.070704f
C522 XA20/CPO D<6> 0.062543f
C523 AVDD XA0/CP0 0.056802f
C524 XA4/CEO XA5/CEO 0.431792f
C525 VREF XA4/EN 0.153675f
C526 SARN XA20/XA3/N1 0.052572f
C527 VREF D<7> 0.08346f
C528 XA0/XA4/A D<8> 0.064665f
C529 XA20/CNO XA3/XA4/A 0.286129f
C530 EN XA2/XA4/A 0.088464f
C531 EN XA5/XA2/A 0.11418f
C532 XA20/CNO D<2> 0.06424f
C533 XA20/CNO XA2/CN1 0.191319f
C534 XA7/CN0 D<3> 0.155005f
C535 XA2/CN0 D<2> 0.072968f
C536 XA2/CN0 XA2/CN1 0.582357f
C537 XA7/EN XA7/XA1/XA1/MP3/G 0.095485f
C538 XA2/EN D<7> 0.084621f
C539 XA3/EN XA3/CN1 0.231584f
C540 XA0/CP0 D<8> 0.113231f
C541 CK_SAMPLE D<4> 0.100705f
C542 VREF D<1> 0.08346f
C543 XA0/XA1/XA2/Y XA20/CPO 0.069784f
C544 XA5/CN0 D<3> 1.413926f
C545 XA2/CN1 XA3/CP0 0.065837f
C546 XA3/EN D<5> 0.063821f
C547 XA7/EN D<1> 0.071215f
C548 AVDD XA1/CEO 0.346648f
C549 XA20/CPO XA6/CN0 0.064431f
C550 XA2/CEO XA3/XA11/A 0.06726f
C551 D<4> XA1/CN0 0.070487f
C552 D<7> XA0/CP0 1.030587f
C553 VREF XA3/EN 0.153675f
C554 XA3/CN0 D<2> 0.069299f
C555 XA2/CN1 XA3/CN0 0.069604f
C556 CK_SAMPLE XA1/CN0 0.071155f
C557 XA2/CEO VREF 0.367402f
C558 XA20/CPO XA2/CP0 0.060601f
C559 XA3/CEO XA3/XA11/A 0.126482f
C560 XA20/CNO D<3> 0.064471f
C561 XA2/CN0 D<3> 0.269469f
C562 XA1/CP0 XA1/CN0 3.110844f
C563 XA8/XA9/MN1/a_324_334# AVSS 0.360976f
C564 XA8/XA9/MN0/a_324_n18# AVSS 0.359088f
C565 XA8/XA9/A AVSS 1.251534f
C566 DONE AVSS 0.857355f
C567 XA8/XA7/MN0/a_324_n18# AVSS 0.359306f
C568 XA8/XA8/MN0/a_324_n18# AVSS 0.360976f
C569 XA8/XA9/B AVSS 1.146132f
C570 XA8/XA6/MN0/a_324_n18# AVSS 0.360779f
C571 XA8/XA4/A AVSS 2.617843f
C572 XA8/XA4/MN0/a_324_n18# AVSS 0.360976f
C573 XA8/CP0 AVSS 2.410423f
C574 XA8/CN0 AVSS 0.310902f
C575 XA8/XA5/MN0/a_324_n18# AVSS 0.360976f
C576 XA8/CN1 AVSS 2.439039f
C577 D<0> AVSS 0.416402f
C578 XA8/XA3/MN0/a_324_n18# AVSS 0.360976f
C579 XA8/XA2/A AVSS 2.029939f
C580 XA8/XA2/MN0/a_324_n18# AVSS 0.359554f
C581 XA8/XA1/XA5/MN0/a_324_n18# AVSS 0.359602f
C582 XA8/XA1/XA4/MN0/a_324_n18# AVSS 0.360806f
C583 XA8/XA1/XA2/MN0/a_324_n18# AVSS 0.360976f
C584 XA8/XA1/XA2/Y AVSS 1.056312f
C585 XA8/XA1/XA1/MN3/a_324_n18# AVSS 0.355765f
C586 XA8/XA1/XA1/MN2/a_324_n18# AVSS 0.355856f
C587 XA8/XA1/XA1/MN1/a_324_n18# AVSS 0.355616f
C588 XA8/XA1/XA1/MP3/G AVSS 0.828529f
C589 XA8/XA1/XA1/MN2/S AVSS 0.200627f
C590 XA8/XA1/XA1/MN0/a_324_n18# AVSS 0.361067f
C591 XA8/ENO AVSS 1.730991f
C592 XA8/XA1/XA0/MN1/a_324_n18# AVSS 0.422745f
C593 XA8/XA1/XA0/MP1/a_216_n18# AVSS 0.091271f
C594 XA8/XA13/MN1/a_324_334# AVSS 0.436861f
C595 XA8/XA13/MP1/a_216_334# AVSS 0.098348f
C596 XA8/XA12/MN0/a_324_n18# AVSS 0.361337f
C597 XA8/XA13/MN1/a_324_n18# AVSS 0.361858f
C598 XA8/XA12/A AVSS 0.761772f
C599 XA8/XA11/MN0/a_324_n18# AVSS 0.360976f
C600 XA7/CEO AVSS 1.549428f
C601 XA8/XA11/A AVSS 0.665842f
C602 XA8/XA9/Y AVSS 0.720752f
C603 XA7/XA9/MN1/a_324_334# AVSS 0.360976f
C604 XA7/XA9/MN0/a_324_n18# AVSS 0.360859f
C605 XA7/XA9/A AVSS 1.253304f
C606 XA7/DONE AVSS 0.085638f
C607 XA7/XA7/MN0/a_324_n18# AVSS 0.360797f
C608 XA7/XA8/MN0/a_324_n18# AVSS 0.360976f
C609 XA7/XA9/B AVSS 1.158973f
C610 XA7/XA6/MN0/a_324_n18# AVSS 0.360724f
C611 XA7/XA4/A AVSS 2.58573f
C612 XA7/XA4/MN0/a_324_n18# AVSS 0.360976f
C613 XA7/CP0 AVSS 2.408835f
C614 XA7/CN0 AVSS 4.433667f
C615 XA7/XA5/MN0/a_324_n18# AVSS 0.360976f
C616 XA7/CN1 AVSS 2.42055f
C617 D<1> AVSS 7.212773f
C618 XA7/XA3/MN0/a_324_n18# AVSS 0.360976f
C619 XA7/XA2/A AVSS 2.012003f
C620 XA7/XA2/MN0/a_324_n18# AVSS 0.359675f
C621 XA7/XA1/XA5/MN0/a_324_n18# AVSS 0.359153f
C622 XA7/XA1/XA4/MN0/a_324_n18# AVSS 0.360841f
C623 XA7/XA1/XA2/MN0/a_324_n18# AVSS 0.360976f
C624 XA7/XA1/XA2/Y AVSS 1.050594f
C625 XA7/XA1/XA1/MN3/a_324_n18# AVSS 0.355765f
C626 XA7/XA1/XA1/MN2/a_324_n18# AVSS 0.353808f
C627 XA7/XA1/XA1/MN1/a_324_n18# AVSS 0.354098f
C628 XA7/XA1/XA1/MP3/G AVSS 0.805069f
C629 XA7/XA1/XA1/MN2/S AVSS 0.168617f
C630 XA7/XA1/XA1/MN0/a_324_n18# AVSS 0.358813f
C631 XA8/EN AVSS 4.2973f
C632 XA7/XA1/XA0/MN1/a_324_n18# AVSS 0.422745f
C633 XA7/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C634 XA7/XA13/MN1/a_324_334# AVSS 0.436861f
C635 XA7/XA13/MP1/a_216_334# AVSS 0.098348f
C636 XA7/XA12/MN0/a_324_n18# AVSS 0.361051f
C637 XA7/XA13/MN1/a_324_n18# AVSS 0.361891f
C638 XA7/XA12/A AVSS 0.719596f
C639 XA7/XA11/MN0/a_324_n18# AVSS 0.360633f
C640 XA6/CEO AVSS 1.369495f
C641 XA7/XA11/A AVSS 0.657884f
C642 XA7/XA9/Y AVSS 0.720752f
C643 XA6/XA9/MN1/a_324_334# AVSS 0.360976f
C644 XA6/XA9/MN0/a_324_n18# AVSS 0.360859f
C645 XA6/XA9/A AVSS 1.253304f
C646 XA6/DONE AVSS 0.085638f
C647 XA6/XA7/MN0/a_324_n18# AVSS 0.360797f
C648 XA6/XA8/MN0/a_324_n18# AVSS 0.360976f
C649 XA6/XA9/B AVSS 1.159109f
C650 XA6/XA6/MN0/a_324_n18# AVSS 0.360724f
C651 XA6/XA4/A AVSS 2.586998f
C652 XA6/XA4/MN0/a_324_n18# AVSS 0.360976f
C653 XA6/CP0 AVSS 2.408736f
C654 XA6/CN0 AVSS 3.681778f
C655 XA6/XA5/MN0/a_324_n18# AVSS 0.360976f
C656 XA6/CN1 AVSS 2.419203f
C657 D<2> AVSS 5.82271f
C658 XA6/XA3/MN0/a_324_n18# AVSS 0.360976f
C659 XA6/XA2/A AVSS 2.011646f
C660 XA6/XA2/MN0/a_324_n18# AVSS 0.359675f
C661 XA6/XA1/XA5/MN0/a_324_n18# AVSS 0.359681f
C662 XA6/XA1/XA4/MN0/a_324_n18# AVSS 0.360841f
C663 XA6/XA1/XA2/MN0/a_324_n18# AVSS 0.360976f
C664 XA6/XA1/XA2/Y AVSS 1.051535f
C665 XA6/XA1/XA1/MN3/a_324_n18# AVSS 0.355765f
C666 XA6/XA1/XA1/MN2/a_324_n18# AVSS 0.355856f
C667 XA6/XA1/XA1/MN1/a_324_n18# AVSS 0.355616f
C668 XA6/XA1/XA1/MP3/G AVSS 0.818898f
C669 XA6/XA1/XA1/MN2/S AVSS 0.192661f
C670 XA6/XA1/XA1/MN0/a_324_n18# AVSS 0.361067f
C671 XA7/EN AVSS 4.111737f
C672 XA6/XA1/XA0/MN1/a_324_n18# AVSS 0.422745f
C673 XA6/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C674 XA6/XA13/MN1/a_324_334# AVSS 0.436861f
C675 XA6/XA13/MP1/a_216_334# AVSS 0.098348f
C676 XA6/XA12/MN0/a_324_n18# AVSS 0.361337f
C677 XA6/XA13/MN1/a_324_n18# AVSS 0.361858f
C678 XA6/XA12/A AVSS 0.761858f
C679 XA6/XA11/MN0/a_324_n18# AVSS 0.360976f
C680 XA5/CEO AVSS 1.548527f
C681 XA6/XA11/A AVSS 0.665857f
C682 XA6/XA9/Y AVSS 0.720752f
C683 XA5/XA9/MN1/a_324_334# AVSS 0.360976f
C684 XA5/XA9/MN0/a_324_n18# AVSS 0.360859f
C685 XA5/XA9/A AVSS 1.253304f
C686 XA5/DONE AVSS 0.085638f
C687 XA5/XA7/MN0/a_324_n18# AVSS 0.360797f
C688 XA5/XA8/MN0/a_324_n18# AVSS 0.360976f
C689 XA5/XA9/B AVSS 1.158973f
C690 XA5/XA6/MN0/a_324_n18# AVSS 0.360724f
C691 XA5/XA4/A AVSS 2.58573f
C692 XA5/XA4/MN0/a_324_n18# AVSS 0.360976f
C693 XA5/CP0 AVSS 2.408835f
C694 XA5/CN0 AVSS 2.651166f
C695 XA5/XA5/MN0/a_324_n18# AVSS 0.360976f
C696 XA5/CN1 AVSS 2.42055f
C697 D<3> AVSS 4.724081f
C698 XA5/XA3/MN0/a_324_n18# AVSS 0.360976f
C699 XA5/XA2/A AVSS 2.012003f
C700 XA5/XA2/MN0/a_324_n18# AVSS 0.359675f
C701 XA5/XA1/XA5/MN0/a_324_n18# AVSS 0.359153f
C702 XA5/XA1/XA4/MN0/a_324_n18# AVSS 0.360841f
C703 XA5/XA1/XA2/MN0/a_324_n18# AVSS 0.360976f
C704 XA5/XA1/XA2/Y AVSS 1.050594f
C705 XA5/XA1/XA1/MN3/a_324_n18# AVSS 0.355765f
C706 XA5/XA1/XA1/MN2/a_324_n18# AVSS 0.353808f
C707 XA5/XA1/XA1/MN1/a_324_n18# AVSS 0.354098f
C708 XA5/XA1/XA1/MP3/G AVSS 0.805069f
C709 XA5/XA1/XA1/MN2/S AVSS 0.168617f
C710 XA5/XA1/XA1/MN0/a_324_n18# AVSS 0.358813f
C711 XA6/EN AVSS 4.241973f
C712 XA5/XA1/XA0/MN1/a_324_n18# AVSS 0.422745f
C713 XA5/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C714 XA5/XA13/MN1/a_324_334# AVSS 0.436861f
C715 XA5/XA13/MP1/a_216_334# AVSS 0.098348f
C716 XA5/XA12/MN0/a_324_n18# AVSS 0.361051f
C717 XA5/XA13/MN1/a_324_n18# AVSS 0.361891f
C718 XA5/XA12/A AVSS 0.719596f
C719 XA5/XA11/MN0/a_324_n18# AVSS 0.360633f
C720 XA4/CEO AVSS 1.369495f
C721 XA5/XA11/A AVSS 0.657884f
C722 XA5/XA9/Y AVSS 0.720752f
C723 XA4/XA9/MN1/a_324_334# AVSS 0.360976f
C724 XA4/XA9/MN0/a_324_n18# AVSS 0.360859f
C725 XA4/XA9/A AVSS 1.253304f
C726 XA4/DONE AVSS 0.085638f
C727 XA4/XA7/MN0/a_324_n18# AVSS 0.360797f
C728 XA4/XA8/MN0/a_324_n18# AVSS 0.360976f
C729 XA4/XA9/B AVSS 1.159109f
C730 XA4/XA6/MN0/a_324_n18# AVSS 0.360724f
C731 XA4/XA4/A AVSS 2.584042f
C732 XA4/XA4/MN0/a_324_n18# AVSS 0.360976f
C733 XA4/CP0 AVSS 2.408736f
C734 XA4/CN0 AVSS 3.172689f
C735 XA4/XA5/MN0/a_324_n18# AVSS 0.360976f
C736 XA4/CN1 AVSS 2.418961f
C737 D<4> AVSS 4.69694f
C738 XA4/XA3/MN0/a_324_n18# AVSS 0.360407f
C739 XA4/XA2/A AVSS 2.006699f
C740 XA4/XA2/MN0/a_324_n18# AVSS 0.359106f
C741 XA4/XA1/XA5/MN0/a_324_n18# AVSS 0.359112f
C742 XA4/XA1/XA4/MN0/a_324_n18# AVSS 0.360272f
C743 XA4/XA1/XA2/MN0/a_324_n18# AVSS 0.360407f
C744 XA4/XA1/XA2/Y AVSS 1.048631f
C745 XA4/XA1/XA1/MN3/a_324_n18# AVSS 0.355196f
C746 XA4/XA1/XA1/MN2/a_324_n18# AVSS 0.355196f
C747 XA4/XA1/XA1/MN1/a_324_n18# AVSS 0.355019f
C748 XA4/XA1/XA1/MP3/G AVSS 0.817852f
C749 XA4/XA1/XA1/MN2/S AVSS 0.192661f
C750 XA4/XA1/XA1/MN0/a_324_n18# AVSS 0.360407f
C751 XA5/EN AVSS 4.122032f
C752 XA4/XA1/XA0/MN1/a_324_n18# AVSS 0.422415f
C753 XA4/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C754 XA4/XA13/MN1/a_324_334# AVSS 0.436861f
C755 XA4/XA13/MP1/a_216_334# AVSS 0.098348f
C756 XA4/XA12/MN0/a_324_n18# AVSS 0.361337f
C757 XA4/XA13/MN1/a_324_n18# AVSS 0.361858f
C758 XA4/XA12/A AVSS 0.761858f
C759 XA4/XA11/MN0/a_324_n18# AVSS 0.360976f
C760 XA3/CEO AVSS 1.548528f
C761 XA4/XA11/A AVSS 0.665857f
C762 XA4/XA9/Y AVSS 0.720752f
C763 XA3/XA9/MN1/a_324_334# AVSS 0.360976f
C764 XA3/XA9/MN0/a_324_n18# AVSS 0.360859f
C765 XA3/XA9/A AVSS 1.253304f
C766 XA3/DONE AVSS 0.085638f
C767 XA3/XA7/MN0/a_324_n18# AVSS 0.360797f
C768 XA3/XA8/MN0/a_324_n18# AVSS 0.360976f
C769 XA3/XA9/B AVSS 1.158973f
C770 XA3/XA6/MN0/a_324_n18# AVSS 0.360724f
C771 XA3/XA4/A AVSS 2.582657f
C772 XA3/XA4/MN0/a_324_n18# AVSS 0.360976f
C773 XA3/CP0 AVSS 4.891468f
C774 XA3/CN0 AVSS 3.451131f
C775 XA3/XA5/MN0/a_324_n18# AVSS 0.360976f
C776 XA3/CN1 AVSS 7.759504f
C777 D<5> AVSS 6.193985f
C778 XA3/XA3/MN0/a_324_n18# AVSS 0.359315f
C779 XA3/XA2/A AVSS 1.990744f
C780 XA3/XA2/MN0/a_324_n18# AVSS 0.358014f
C781 XA3/XA1/XA5/MN0/a_324_n18# AVSS 0.357579f
C782 XA3/XA1/XA4/MN0/a_324_n18# AVSS 0.35918f
C783 XA3/XA1/XA2/MN0/a_324_n18# AVSS 0.359315f
C784 XA3/XA1/XA2/Y AVSS 1.041199f
C785 XA3/XA1/XA1/MN3/a_324_n18# AVSS 0.354104f
C786 XA3/XA1/XA1/MN2/a_324_n18# AVSS 0.352056f
C787 XA3/XA1/XA1/MN1/a_324_n18# AVSS 0.352346f
C788 XA3/XA1/XA1/MP3/G AVSS 0.800747f
C789 XA3/XA1/XA1/MN2/S AVSS 0.168617f
C790 XA3/XA1/XA1/MN0/a_324_n18# AVSS 0.357093f
C791 XA4/EN AVSS 4.2646f
C792 XA3/XA1/XA0/MN1/a_324_n18# AVSS 0.421869f
C793 XA3/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C794 XA3/XA13/MN1/a_324_334# AVSS 0.436861f
C795 XA3/XA13/MP1/a_216_334# AVSS 0.098348f
C796 XA3/XA12/MN0/a_324_n18# AVSS 0.361051f
C797 XA3/XA13/MN1/a_324_n18# AVSS 0.361891f
C798 XA3/XA12/A AVSS 0.719596f
C799 XA3/XA11/MN0/a_324_n18# AVSS 0.360633f
C800 XA2/CEO AVSS 1.368725f
C801 XA3/XA11/A AVSS 0.657884f
C802 XA3/XA9/Y AVSS 0.720752f
C803 XA2/XA9/MN1/a_324_334# AVSS 0.360976f
C804 XA2/XA9/MN0/a_324_n18# AVSS 0.360859f
C805 XA2/XA9/A AVSS 1.253304f
C806 XA2/DONE AVSS 0.085638f
C807 XA2/XA7/MN0/a_324_n18# AVSS 0.360797f
C808 XA2/XA8/MN0/a_324_n18# AVSS 0.360976f
C809 XA2/XA9/B AVSS 1.159109f
C810 XA2/XA6/MN0/a_324_n18# AVSS 0.360724f
C811 XA2/XA4/A AVSS 2.583863f
C812 XA2/XA4/MN0/a_324_n18# AVSS 0.360976f
C813 XA2/CP0 AVSS 4.847463f
C814 XA2/CN0 AVSS 3.206913f
C815 XA2/XA5/MN0/a_324_n18# AVSS 0.360976f
C816 XA2/CN1 AVSS 6.009428f
C817 D<6> AVSS 5.15921f
C818 XA2/XA3/MN0/a_324_n18# AVSS 0.359924f
C819 XA2/XA2/A AVSS 2.00081f
C820 XA2/XA2/MN0/a_324_n18# AVSS 0.358622f
C821 XA2/XA1/XA5/MN0/a_324_n18# AVSS 0.358629f
C822 XA2/XA1/XA4/MN0/a_324_n18# AVSS 0.359789f
C823 XA2/XA1/XA2/MN0/a_324_n18# AVSS 0.359924f
C824 XA2/XA1/XA2/Y AVSS 1.046445f
C825 XA2/XA1/XA1/MN3/a_324_n18# AVSS 0.354713f
C826 XA2/XA1/XA1/MN2/a_324_n18# AVSS 0.354713f
C827 XA2/XA1/XA1/MN1/a_324_n18# AVSS 0.354713f
C828 XA2/XA1/XA1/MP3/G AVSS 0.816518f
C829 XA2/XA1/XA1/MN2/S AVSS 0.192661f
C830 XA2/XA1/XA1/MN0/a_324_n18# AVSS 0.359924f
C831 XA3/EN AVSS 4.173967f
C832 XA2/XA1/XA0/MN1/a_324_n18# AVSS 0.422173f
C833 XA2/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C834 XA2/XA13/MN1/a_324_334# AVSS 0.436861f
C835 XA2/XA13/MP1/a_216_334# AVSS 0.098348f
C836 XA2/XA12/MN0/a_324_n18# AVSS 0.361337f
C837 XA2/XA13/MN1/a_324_n18# AVSS 0.361858f
C838 XA2/XA12/A AVSS 0.761858f
C839 XA2/XA11/MN0/a_324_n18# AVSS 0.360976f
C840 XA1/CEO AVSS 1.548527f
C841 XA2/XA11/A AVSS 0.665857f
C842 XA2/XA9/Y AVSS 0.720752f
C843 XB2/XA7/MN1/a_324_n18# AVSS 0.359583f
C844 XB2/XA5b/MN1/a_324_n18# AVSS 0.436157f
C845 XB2/XA0/MN0/a_324_n18# AVSS 0.359945f
C846 XB2/XA5b/MP1/a_216_n18# AVSS 0.098348f
C847 XB2/XA1/Y AVSS 0.690192f
C848 XB2/XA4/MN1/a_324_334# AVSS 0.359583f
C849 XB2/XA4/MN0/a_324_n18# AVSS 0.359583f
C850 XB2/XA5/MN1/a_324_334# AVSS 0.422f
C851 XB2/XA5/MP1/a_216_334# AVSS 0.091271f
C852 XB2/XA3/B AVSS 55.474865f
C853 XB2/XA3/MP0/S AVSS 0.744149f
C854 XB2/XA7/MN1/a_324_334# AVSS 0.359583f
C855 XB2/XA5/MN1/a_324_n18# AVSS 0.360407f
C856 XB2/XA2/MP0/G AVSS 0.708335f
C857 XB2/XA1/MP0/G AVSS 0.788614f
C858 XB2/XA3/MN0/a_324_n18# AVSS 0.359855f
C859 XB2/CKN AVSS 1.785976f
C860 XB2/M8/a_324_n18# AVSS 0.356455f
C861 XB2/M8/a_324_334# AVSS 0.421527f
C862 XB2/M7/a_324_n18# AVSS 0.356455f
C863 XB2/XA4/GNG AVSS 54.21507f
C864 XB2/M6/a_324_n18# AVSS 0.356455f
C865 XB2/M3/a_324_n18# AVSS 0.356755f
C866 XB2/M4/a_324_n18# AVSS 0.35654f
C867 XB2/M5/a_324_n18# AVSS 0.356434f
C868 XB2/M2/a_324_n18# AVSS 0.357028f
C869 XB2/M4/G AVSS 2.47803f
C870 SAR_IN AVSS 1.183928f
C871 XB2/M1/a_324_n18# AVSS 0.429021f
C872 XA1/XA9/MN1/a_324_334# AVSS 0.360976f
C873 XA1/XA9/MN0/a_324_n18# AVSS 0.360859f
C874 XA1/XA9/A AVSS 1.253304f
C875 XA1/DONE AVSS 0.085638f
C876 XA1/XA7/MN0/a_324_n18# AVSS 0.360797f
C877 XA1/XA8/MN0/a_324_n18# AVSS 0.360976f
C878 XA1/XA9/B AVSS 1.158973f
C879 XA1/XA6/MN0/a_324_n18# AVSS 0.360724f
C880 XA1/XA4/A AVSS 2.582657f
C881 XA1/XA4/MN0/a_324_n18# AVSS 0.360976f
C882 XA1/CP0 AVSS 8.128386f
C883 XA1/XA5/MN0/a_324_n18# AVSS 0.360976f
C884 XA1/CN1 AVSS 8.016429f
C885 XA1/XA3/MN0/a_324_n18# AVSS 0.359047f
C886 VREF AVSS 34.767807f
C887 XA1/XA2/A AVSS 1.987538f
C888 XA1/XA2/MN0/a_324_n18# AVSS 0.357746f
C889 XA1/XA1/XA5/MN0/a_324_n18# AVSS 0.357311f
C890 XA1/XA1/XA4/MN0/a_324_n18# AVSS 0.358912f
C891 XA1/XA1/XA2/MN0/a_324_n18# AVSS 0.359047f
C892 XA1/XA1/XA2/Y AVSS 1.039978f
C893 XA1/XA1/XA1/MN3/a_324_n18# AVSS 0.353836f
C894 XA1/XA1/XA1/MN2/a_324_n18# AVSS 0.351788f
C895 XA1/XA1/XA1/MN1/a_324_n18# AVSS 0.352078f
C896 XA1/XA1/XA1/MP3/G AVSS 0.800137f
C897 XA1/XA1/XA1/MN2/S AVSS 0.168617f
C898 XA1/XA1/XA1/MN0/a_324_n18# AVSS 0.356825f
C899 XA2/EN AVSS 4.229634f
C900 XA1/XA1/XA0/MN1/a_324_n18# AVSS 0.421735f
C901 XA1/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C902 XA1/XA13/MN1/a_324_334# AVSS 0.436861f
C903 XA1/XA13/MP1/a_216_334# AVSS 0.098348f
C904 XA1/XA12/MN0/a_324_n18# AVSS 0.361051f
C905 XA1/XA13/MN1/a_324_n18# AVSS 0.361891f
C906 XA1/XA12/A AVSS 0.719596f
C907 XA1/XA11/MN0/a_324_n18# AVSS 0.360633f
C908 XA0/CEO AVSS 1.367197f
C909 XA1/XA11/A AVSS 0.657884f
C910 XA1/XA9/Y AVSS 0.720752f
C911 XA0/XA9/MN1/a_324_334# AVSS 0.361065f
C912 XA0/XA9/MN0/a_324_n18# AVSS 0.360745f
C913 XA0/XA9/A AVSS 1.251784f
C914 XA0/DONE AVSS 0.085638f
C915 XA0/XA7/MN0/a_324_n18# AVSS 0.36065f
C916 XA0/XA8/MN0/a_324_n18# AVSS 0.36083f
C917 XA0/XA9/B AVSS 1.20293f
C918 CK_SAMPLE AVSS 20.221697f
C919 XA0/XA6/MN0/a_324_n18# AVSS 0.360781f
C920 XA0/XA4/A AVSS 2.658212f
C921 XA0/XA4/MN0/a_324_n18# AVSS 0.36083f
C922 XA0/XA5/MN0/a_324_n18# AVSS 0.361065f
C923 XA0/XA3/MN0/a_324_n18# AVSS 0.360346f
C924 XA0/XA2/A AVSS 2.00376f
C925 XA0/XA2/MN0/a_324_n18# AVSS 0.359045f
C926 XA0/XA1/XA5/MN0/a_324_n18# AVSS 0.35872f
C927 EN AVSS 7.481703f
C928 XA0/XA1/XA4/MN0/a_324_n18# AVSS 0.35988f
C929 XA0/XA1/XA2/MN0/a_324_n18# AVSS 0.360015f
C930 XA0/XA1/XA2/Y AVSS 1.046893f
C931 XA0/XA1/XA1/MN3/a_324_n18# AVSS 0.354804f
C932 XA20/CPO AVSS 14.364732f
C933 XA0/XA1/XA1/MN2/a_324_n18# AVSS 0.354804f
C934 XA20/CNO AVSS 15.685797f
C935 XA0/XA1/XA1/MN1/a_324_n18# AVSS 0.354804f
C936 XA0/XA1/XA1/MP3/G AVSS 0.817052f
C937 XA0/XA1/XA1/MN2/S AVSS 0.192661f
C938 XA0/XA1/XA1/MN0/a_324_n18# AVSS 0.36064f
C939 XA1/EN AVSS 4.171568f
C940 XA0/XA1/XA0/MN1/a_324_n18# AVSS 0.42289f
C941 AVDD AVSS 0.582587p
C942 XA0/XA1/XA0/MP1/a_216_n18# AVSS 0.091111f
C943 XA0/XA13/MN1/a_324_334# AVSS 0.436917f
C944 XA0/XA13/MP1/a_216_334# AVSS 0.098348f
C945 XA0/XA12/MN0/a_324_n18# AVSS 0.361426f
C946 XA0/XA13/MN1/a_324_n18# AVSS 0.361914f
C947 XA0/XA12/A AVSS 0.760999f
C948 XA0/XA11/MN0/a_324_n18# AVSS 0.361065f
C949 XA0/XA11/A AVSS 0.665137f
C950 XA0/XA9/Y AVSS 0.719968f
C951 XB1/XA7/MN1/a_324_n18# AVSS 0.359583f
C952 XB1/XA5b/MN1/a_324_n18# AVSS 0.436157f
C953 XB1/XA0/MN0/a_324_n18# AVSS 0.359977f
C954 XB1/XA5b/MP1/a_216_n18# AVSS 0.098348f
C955 XB1/XA1/Y AVSS 0.690192f
C956 XB1/XA4/MN1/a_324_334# AVSS 0.359583f
C957 XB1/XA4/MN0/a_324_n18# AVSS 0.359583f
C958 XB1/XA5/MN1/a_324_334# AVSS 0.422f
C959 XB1/XA5/MP1/a_216_334# AVSS 0.091271f
C960 XB1/XA3/B AVSS 55.47486f
C961 XB1/XA3/MP0/S AVSS 0.744194f
C962 XB1/XA7/MN1/a_324_334# AVSS 0.359583f
C963 XB1/XA5/MN1/a_324_n18# AVSS 0.360407f
C964 XB1/XA2/MP0/G AVSS 0.708335f
C965 XB1/XA1/MP0/G AVSS 0.788614f
C966 XB1/XA3/MN0/a_324_n18# AVSS 0.359873f
C967 CK_SAMPLE_BSSW AVSS 4.64133f
C968 XB1/CKN AVSS 1.786059f
C969 XB1/M8/a_324_n18# AVSS 0.356455f
C970 XB1/M8/a_324_334# AVSS 0.421527f
C971 XB1/M7/a_324_n18# AVSS 0.356455f
C972 XA0/CEIN AVSS 29.52815f
C973 XB1/XA4/GNG AVSS 54.21506f
C974 XB1/M6/a_324_n18# AVSS 0.356455f
C975 XB1/M3/a_324_n18# AVSS 0.356755f
C976 XB1/M4/a_324_n18# AVSS 0.35654f
C977 XB1/M5/a_324_n18# AVSS 0.356434f
C978 XB1/M2/a_324_n18# AVSS 0.357028f
C979 SARP AVSS 47.616425f
C980 XB1/M4/G AVSS 2.475204f
C981 SAR_IP AVSS 1.183778f
C982 XB1/M1/a_324_n18# AVSS 0.429021f
C983 XA20/XA9/MN0/a_324_n18# AVSS 0.360499f
C984 XA20/XA3/CO AVSS 2.696206f
C985 XA20/XA2/MN6/a_324_334# AVSS 0.360239f
C986 XA20/XA3a/A AVSS 2.538063f
C987 XA20/XA3/MN0/a_324_n18# AVSS 0.360499f
C988 XA20/XA3a/MN0/a_324_n18# AVSS 0.360319f
C989 XA20/XA4/MN0/a_324_n18# AVSS 0.360499f
C990 XA20/XA4/MP0/S AVSS 0.397005f
C991 SARN AVSS 48.72758f
C992 XA20/XA3/N2 AVSS 0.234927f
C993 XA20/XA9/Y AVSS 3.177331f
C994 XA20/XA2/N2 AVSS 0.234927f
C995 XA20/XA2/MN0/a_324_n18# AVSS 0.360499f
C996 XA20/XA3/N1 AVSS 0.904779f
C997 XA20/XA1/MN0/a_324_n18# AVSS 0.359764f
C998 XA20/XA1/MP0/S AVSS 0.397011f
C999 XA20/XA9/A AVSS 3.901928f
C1000 XA20/XA0/MN1/a_324_n18# AVSS 0.422452f
C1001 XA20/XA0/MP1/a_216_n18# AVSS 0.091271f
C1002 XA20/XA13/MN1/a_324_334# AVSS 0.433288f
C1003 XA20/XA13/MP1/a_216_334# AVSS 0.092623f
C1004 XA20/XA13/MN1/a_324_n18# AVSS 0.361124f
C1005 XA8/CEO AVSS 1.013552f
C1006 XA20/XA12/MN0/a_324_n18# AVSS 0.361124f
C1007 XA20/XA11/MN0/a_324_n18# AVSS 0.361068f
C1008 XA20/XA9/MN0/a_324_334# AVSS 0.36083f
C1009 XA20/XA12/Y AVSS 0.624428f
C1010 XA20/XA11/Y AVSS 0.761175f
C1011 XA0/CN0 AVSS 10.220659f
C1012 XA1/CN0 AVSS 6.575425f
C1013 D<8> AVSS 11.982146f
C1014 XDAC2/XC32a<0>/XRES16/B AVSS 4.882681f
C1015 XDAC2/XC32a<0>/XRES8/B AVSS 4.160893f
C1016 XDAC2/XC32a<0>/XRES4/B AVSS 3.745652f
C1017 XDAC2/XC32a<0>/XRES1B/B AVSS 3.315972f
C1018 XDAC2/XC32a<0>/XRES1A/B AVSS 1.751315f
C1019 XDAC2/XC32a<0>/XRES2/B AVSS 3.488831f
C1020 XDAC2/XC128a<1>/XRES16/B AVSS 4.882681f
C1021 XDAC2/XC128a<1>/XRES8/B AVSS 4.160893f
C1022 XDAC2/XC128a<1>/XRES4/B AVSS 3.745652f
C1023 XDAC2/XC128a<1>/XRES1B/B AVSS 3.315972f
C1024 XDAC2/XC128a<1>/XRES1A/B AVSS 1.751315f
C1025 XDAC2/XC128a<1>/XRES2/B AVSS 3.488831f
C1026 XDAC2/XC64b<1>/XRES16/B AVSS 4.882681f
C1027 XDAC2/XC64b<1>/XRES8/B AVSS 4.160893f
C1028 XDAC2/XC64b<1>/XRES4/B AVSS 3.745652f
C1029 XDAC2/XC64b<1>/XRES1B/B AVSS 3.315972f
C1030 XDAC2/XC64b<1>/XRES1A/B AVSS 1.751315f
C1031 XDAC2/XC64b<1>/XRES2/B AVSS 3.488831f
C1032 XDAC2/XC1/XRES16/B AVSS 4.882681f
C1033 XDAC2/XC1/XRES8/B AVSS 4.160893f
C1034 XDAC2/XC1/XRES4/B AVSS 3.745652f
C1035 XDAC2/XC1/XRES1B/B AVSS 3.315972f
C1036 XDAC2/XC1/XRES1A/B AVSS 1.751315f
C1037 XDAC2/XC1/XRES2/B AVSS 3.488831f
C1038 XDAC2/XC0/XRES16/B AVSS 4.882681f
C1039 XDAC2/XC0/XRES8/B AVSS 4.160893f
C1040 XDAC2/XC0/XRES4/B AVSS 3.745652f
C1041 XDAC2/XC0/XRES1B/B AVSS 3.315972f
C1042 XDAC2/XC0/XRES1A/B AVSS 1.751315f
C1043 XDAC2/XC0/XRES2/B AVSS 3.488831f
C1044 XDAC2/XC64a<0>/XRES16/B AVSS 4.88268f
C1045 XDAC2/XC64a<0>/XRES8/B AVSS 4.160893f
C1046 XDAC2/XC64a<0>/XRES4/B AVSS 3.745652f
C1047 XDAC2/XC64a<0>/XRES1B/B AVSS 3.315972f
C1048 XDAC2/XC64a<0>/XRES1A/B AVSS 1.751315f
C1049 XDAC2/XC64a<0>/XRES2/B AVSS 3.488831f
C1050 XDAC2/X16ab/XRES16/B AVSS 4.882681f
C1051 XDAC2/X16ab/XRES8/B AVSS 4.160893f
C1052 XDAC2/X16ab/XRES4/B AVSS 3.745652f
C1053 XDAC2/X16ab/XRES1B/B AVSS 3.315972f
C1054 XDAC2/X16ab/XRES1A/B AVSS 1.751315f
C1055 XDAC2/X16ab/XRES2/B AVSS 3.488831f
C1056 XDAC2/XC128b<2>/XRES16/B AVSS 4.882681f
C1057 XDAC2/XC128b<2>/XRES8/B AVSS 4.160893f
C1058 XDAC2/XC128b<2>/XRES4/B AVSS 3.745652f
C1059 XDAC2/XC128b<2>/XRES1B/B AVSS 3.315972f
C1060 XDAC2/XC128b<2>/XRES1A/B AVSS 1.751315f
C1061 XDAC2/XC128b<2>/XRES2/B AVSS 3.488831f
C1062 XA0/CP0 AVSS 11.743839f
C1063 XA0/CP1 AVSS 10.640906f
C1064 D<7> AVSS 6.648342f
C1065 XDAC1/XC32a<0>/XRES16/B AVSS 4.882681f
C1066 XDAC1/XC32a<0>/XRES8/B AVSS 4.160893f
C1067 XDAC1/XC32a<0>/XRES4/B AVSS 3.745652f
C1068 XDAC1/XC32a<0>/XRES1B/B AVSS 3.315972f
C1069 XDAC1/XC32a<0>/XRES1A/B AVSS 1.751315f
C1070 XDAC1/XC32a<0>/XRES2/B AVSS 3.488831f
C1071 XDAC1/XC128a<1>/XRES16/B AVSS 4.882681f
C1072 XDAC1/XC128a<1>/XRES8/B AVSS 4.160893f
C1073 XDAC1/XC128a<1>/XRES4/B AVSS 3.745652f
C1074 XDAC1/XC128a<1>/XRES1B/B AVSS 3.315972f
C1075 XDAC1/XC128a<1>/XRES1A/B AVSS 1.751315f
C1076 XDAC1/XC128a<1>/XRES2/B AVSS 3.488831f
C1077 XDAC1/XC64b<1>/XRES16/B AVSS 4.882681f
C1078 XDAC1/XC64b<1>/XRES8/B AVSS 4.160893f
C1079 XDAC1/XC64b<1>/XRES4/B AVSS 3.745652f
C1080 XDAC1/XC64b<1>/XRES1B/B AVSS 3.315972f
C1081 XDAC1/XC64b<1>/XRES1A/B AVSS 1.751315f
C1082 XDAC1/XC64b<1>/XRES2/B AVSS 3.488831f
C1083 XDAC1/XC1/XRES16/B AVSS 4.882681f
C1084 XDAC1/XC1/XRES8/B AVSS 4.160893f
C1085 XDAC1/XC1/XRES4/B AVSS 3.745652f
C1086 XDAC1/XC1/XRES1B/B AVSS 3.315972f
C1087 XDAC1/XC1/XRES1A/B AVSS 1.751315f
C1088 XDAC1/XC1/XRES2/B AVSS 3.488831f
C1089 XDAC1/XC0/XRES16/B AVSS 4.882681f
C1090 XDAC1/XC0/XRES8/B AVSS 4.160893f
C1091 XDAC1/XC0/XRES4/B AVSS 3.745652f
C1092 XDAC1/XC0/XRES1B/B AVSS 3.315972f
C1093 XDAC1/XC0/XRES1A/B AVSS 1.751315f
C1094 XDAC1/XC0/XRES2/B AVSS 3.488831f
C1095 XDAC1/XC64a<0>/XRES16/B AVSS 4.88268f
C1096 XDAC1/XC64a<0>/XRES8/B AVSS 4.160893f
C1097 XDAC1/XC64a<0>/XRES4/B AVSS 3.745652f
C1098 XDAC1/XC64a<0>/XRES1B/B AVSS 3.315972f
C1099 XDAC1/XC64a<0>/XRES1A/B AVSS 1.751315f
C1100 XDAC1/XC64a<0>/XRES2/B AVSS 3.488831f
C1101 XDAC1/X16ab/XRES16/B AVSS 4.882681f
C1102 XDAC1/X16ab/XRES8/B AVSS 4.160893f
C1103 XDAC1/X16ab/XRES4/B AVSS 3.745652f
C1104 XDAC1/X16ab/XRES1B/B AVSS 3.315972f
C1105 XDAC1/X16ab/XRES1A/B AVSS 1.751315f
C1106 XDAC1/X16ab/XRES2/B AVSS 3.488831f
C1107 XDAC1/XC128b<2>/XRES16/B AVSS 4.882681f
C1108 XDAC1/XC128b<2>/XRES8/B AVSS 4.160893f
C1109 XDAC1/XC128b<2>/XRES4/B AVSS 3.745652f
C1110 XDAC1/XC128b<2>/XRES1B/B AVSS 3.315972f
C1111 XDAC1/XC128b<2>/XRES1A/B AVSS 1.751315f
C1112 XDAC1/XC128b<2>/XRES2/B AVSS 3.488831f
.ends

