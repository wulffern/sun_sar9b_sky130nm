magic
tech sky130A
magscale 1 2
timestamp 1708902000
<< checkpaint >>
rect 0 0 2520 704
<< locali >>
rect 830 230 898 298
rect 830 406 898 474
rect 1622 406 1690 474
rect 864 582 1032 650
rect 1032 582 1656 650
rect 1032 582 1100 650
rect 1420 54 1656 122
rect 1420 406 1656 474
rect 1420 54 1488 474
rect 756 406 1764 474
rect 324 318 540 386
rect 1980 494 2196 562
rect 324 494 540 562
rect 324 142 540 210
rect 756 582 972 650
rect 2412 308 2628 396
rect -108 308 108 396
<< poly >>
rect 324 334 2196 370
rect 324 158 2196 194
<< m3 >>
rect 1548 0 1732 704
rect 756 0 940 704
rect 1548 0 1732 704
rect 756 0 940 704
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 176
box 0 176 1260 528
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_PCHDL MP2 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP0 
transform 1 0 1260 0 1 176
box 1260 176 2520 528
use SUNSAR_PCHDL MP1 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 230
box 1548 230 1732 298
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 1548 0 1 230
box 1548 230 1732 298
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 756 0 1 54
box 756 54 940 122
<< labels >>
flabel locali s 324 318 540 386 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 1980 494 2196 562 0 FreeSans 400 0 0 0 CN
port 3 nsew signal bidirectional
flabel locali s 324 494 540 562 0 FreeSans 400 0 0 0 C
port 2 nsew signal bidirectional
flabel locali s 324 142 540 210 0 FreeSans 400 0 0 0 RN
port 4 nsew signal bidirectional
flabel locali s 756 582 972 650 0 FreeSans 400 0 0 0 Y
port 5 nsew signal bidirectional
flabel locali s 2412 308 2628 396 0 FreeSans 400 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -108 308 108 396 0 FreeSans 400 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel m3 s 1548 0 1732 704 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 756 0 940 704 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 704
<< end >>
