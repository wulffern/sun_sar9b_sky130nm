magic
tech sky130B
timestamp 1708692311
<< poly >>
rect 162 79 1098 97
<< locali >>
rect 378 291 828 325
rect 216 247 334 281
rect 1044 247 1162 281
rect 199 71 233 193
rect 300 61 334 247
rect 415 203 882 237
rect 415 115 449 149
rect 811 115 845 149
rect 1128 105 1162 247
rect 990 71 1162 105
rect 300 27 828 61
<< metal3 >>
rect 378 0 470 352
rect 774 149 866 352
rect 912 159 1044 193
rect 912 149 946 159
rect 774 115 946 149
rect 774 0 866 115
use SUNSAR_NCHDL  MN0
timestamp 1708642800
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_NCHDL  MN1
timestamp 1708642800
transform 1 0 0 0 1 88
box -90 -66 630 242
use SUNSAR_NCHDL  MN2
timestamp 1708642800
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNSAR_PCHDL  MP0
timestamp 1708642800
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_PCHDL  MP1_DMY
timestamp 1708642800
transform 1 0 630 0 1 88
box 0 -66 720 242
use SUNSAR_PCHDL  MP2
timestamp 1708642800
transform 1 0 630 0 1 176
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1708642800
transform 1 0 774 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1708642800
transform 1 0 990 0 1 159
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut2
timestamp 1708642800
transform 1 0 774 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut3
timestamp 1708642800
transform 1 0 378 0 1 115
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut4
timestamp 1708642800
transform 1 0 378 0 1 115
box 0 0 92 34
<< labels >>
flabel locali s 990 71 1098 105 0 FreeSans 200 0 0 0 C
port 1 nsew signal bidirectional
flabel locali s 774 203 882 237 0 FreeSans 200 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 378 291 486 325 0 FreeSans 200 0 0 0 A
port 2 nsew signal bidirectional
flabel metal3 s 774 0 866 352 0 FreeSans 200 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel metal3 s 378 0 470 352 0 FreeSans 200 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 352
<< end >>
