magic
tech sky130B
magscale 1 2
timestamp 1708383600
<< checkpaint >>
rect -108 0 22680 4224
<< locali >>
rect 20484 1198 20700 1266
rect 20484 494 20700 562
rect 20916 2342 21132 2410
rect 20916 3574 21132 3642
rect 20916 2694 21132 2762
rect 324 1374 540 1442
rect 4500 1374 4716 1442
rect 5364 1374 5580 1442
rect 9540 1374 9756 1442
rect 10404 1374 10620 1442
rect 14580 1374 14796 1442
rect 15444 1374 15660 1442
rect 19620 1374 19836 1442
rect 756 4102 972 4170
rect 4068 4102 4284 4170
rect 5796 4102 6012 4170
rect 9108 4102 9324 4170
rect 10836 4102 11052 4170
rect 14148 4102 14364 4170
rect 15876 4102 16092 4170
rect 19188 4102 19404 4170
rect 324 494 540 562
rect 2412 484 2628 572
rect -108 484 108 572
use SUNSAR_DFRNQNX1_CV XB07 
transform 1 0 0 0 1 0
box 0 0 2520 4224
use SUNSAR_DFRNQNX1_CV XC08 
transform -1 0 5040 0 1 0
box 5040 0 7560 4224
use SUNSAR_DFRNQNX1_CV XD09 
transform 1 0 5040 0 1 0
box 5040 0 7560 4224
use SUNSAR_DFRNQNX1_CV XE10 
transform -1 0 10080 0 1 0
box 10080 0 12600 4224
use SUNSAR_DFRNQNX1_CV XF11 
transform 1 0 10080 0 1 0
box 10080 0 12600 4224
use SUNSAR_DFRNQNX1_CV XG12 
transform -1 0 15120 0 1 0
box 15120 0 17640 4224
use SUNSAR_DFRNQNX1_CV XH13 
transform 1 0 15120 0 1 0
box 15120 0 17640 4224
use SUNSAR_DFRNQNX1_CV XI14 
transform -1 0 20160 0 1 0
box 20160 0 22680 4224
use SUNSAR_TAPCELLB_CV XA1 
transform 1 0 20160 0 1 0
box 20160 0 22680 352
use SUNSAR_IVX1_CV XA2 
transform 1 0 20160 0 1 352
box 20160 352 22680 704
use SUNSAR_IVX1_CV XA3 
transform 1 0 20160 0 1 704
box 20160 704 22680 1056
use SUNSAR_BFX1_CV XA4 
transform 1 0 20160 0 1 1056
box 20160 1056 22680 1584
use SUNSAR_ORX1_CV XA5 
transform 1 0 20160 0 1 1584
box 20160 1584 22680 2464
use SUNSAR_IVX1_CV XA5a 
transform 1 0 20160 0 1 2464
box 20160 2464 22680 2816
use SUNSAR_ANX1_CV XA6 
transform 1 0 20160 0 1 2816
box 20160 2816 22680 3696
<< labels >>
flabel locali s 20484 1198 20700 1266 0 FreeSans 400 0 0 0 CKS
port 1 nsew signal bidirectional
flabel locali s 20484 494 20700 562 0 FreeSans 400 0 0 0 ENABLE
port 2 nsew signal bidirectional
flabel locali s 20916 2342 21132 2410 0 FreeSans 400 0 0 0 CK_SAMPLE
port 3 nsew signal bidirectional
flabel locali s 20916 3574 21132 3642 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 4 nsew signal bidirectional
flabel locali s 20916 2694 21132 2762 0 FreeSans 400 0 0 0 EN
port 5 nsew signal bidirectional
flabel locali s 324 1374 540 1442 0 FreeSans 400 0 0 0 D<7>
port 6 nsew signal bidirectional
flabel locali s 4500 1374 4716 1442 0 FreeSans 400 0 0 0 D<6>
port 7 nsew signal bidirectional
flabel locali s 5364 1374 5580 1442 0 FreeSans 400 0 0 0 D<5>
port 8 nsew signal bidirectional
flabel locali s 9540 1374 9756 1442 0 FreeSans 400 0 0 0 D<4>
port 9 nsew signal bidirectional
flabel locali s 10404 1374 10620 1442 0 FreeSans 400 0 0 0 D<3>
port 10 nsew signal bidirectional
flabel locali s 14580 1374 14796 1442 0 FreeSans 400 0 0 0 D<2>
port 11 nsew signal bidirectional
flabel locali s 15444 1374 15660 1442 0 FreeSans 400 0 0 0 D<1>
port 12 nsew signal bidirectional
flabel locali s 19620 1374 19836 1442 0 FreeSans 400 0 0 0 D<0>
port 13 nsew signal bidirectional
flabel locali s 756 4102 972 4170 0 FreeSans 400 0 0 0 DO<7>
port 14 nsew signal bidirectional
flabel locali s 4068 4102 4284 4170 0 FreeSans 400 0 0 0 DO<6>
port 15 nsew signal bidirectional
flabel locali s 5796 4102 6012 4170 0 FreeSans 400 0 0 0 DO<5>
port 16 nsew signal bidirectional
flabel locali s 9108 4102 9324 4170 0 FreeSans 400 0 0 0 DO<4>
port 17 nsew signal bidirectional
flabel locali s 10836 4102 11052 4170 0 FreeSans 400 0 0 0 DO<3>
port 18 nsew signal bidirectional
flabel locali s 14148 4102 14364 4170 0 FreeSans 400 0 0 0 DO<2>
port 19 nsew signal bidirectional
flabel locali s 15876 4102 16092 4170 0 FreeSans 400 0 0 0 DO<1>
port 20 nsew signal bidirectional
flabel locali s 19188 4102 19404 4170 0 FreeSans 400 0 0 0 DO<0>
port 21 nsew signal bidirectional
flabel locali s 324 494 540 562 0 FreeSans 400 0 0 0 DONE
port 22 nsew signal bidirectional
flabel locali s 2412 484 2628 572 0 FreeSans 400 0 0 0 AVDD
port 23 nsew signal bidirectional
flabel locali s -108 484 108 572 0 FreeSans 400 0 0 0 AVSS
port 24 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -108 22680 0 4224
<< end >>
