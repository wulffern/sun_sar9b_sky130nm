magic
tech sky130B
magscale 1 2
timestamp 1708297200
<< checkpaint >>
rect 0 0 8712 1056
<< m1 >>
rect 108 -44 8676 44
rect 8604 44 8676 132
rect 108 132 8532 220
rect 8604 132 8676 220
rect 108 220 180 308
rect 8604 220 8676 308
rect 108 308 180 396
rect 252 308 8676 396
rect 108 396 180 484
rect 8604 396 8676 484
rect 108 484 8532 572
rect 8604 484 8676 572
rect 108 572 180 660
rect 8604 572 8676 660
rect 108 660 180 748
rect 252 660 8676 748
rect 108 748 180 836
rect 108 836 8676 924
<< m2 >>
rect 108 -44 8676 44
rect 8604 44 8676 132
rect 108 132 8532 220
rect 8604 132 8676 220
rect 108 220 180 308
rect 8604 220 8676 308
rect 108 308 180 396
rect 252 308 8676 396
rect 108 396 180 484
rect 8604 396 8676 484
rect 108 484 8532 572
rect 8604 484 8676 572
rect 108 572 180 660
rect 8604 572 8676 660
rect 108 660 180 748
rect 252 660 8676 748
rect 108 748 180 836
rect 108 836 8676 924
<< locali >>
rect 108 -44 8676 44
rect 8604 44 8676 132
rect 108 132 8532 220
rect 8604 132 8676 220
rect 108 220 180 308
rect 8604 220 8676 308
rect 108 308 180 396
rect 252 308 8676 396
rect 108 396 180 484
rect 8604 396 8676 484
rect 108 484 8532 572
rect 8604 484 8676 572
rect 108 572 180 660
rect 8604 572 8676 660
rect 108 660 180 748
rect 252 660 8676 748
rect 108 748 180 836
rect 108 836 8676 924
<< v1 >>
rect 8316 -35 8388 -26
rect 8316 -26 8388 -17
rect 8316 -17 8388 -8
rect 8316 -8 8388 0
rect 8316 0 8388 8
rect 8316 8 8388 17
rect 8316 17 8388 26
rect 8316 26 8388 35
rect 8388 -35 8460 -26
rect 8388 -26 8460 -17
rect 8388 -17 8460 -8
rect 8388 -8 8460 0
rect 8388 0 8460 8
rect 8388 8 8460 17
rect 8388 17 8460 26
rect 8388 26 8460 35
rect 8460 -35 8532 -26
rect 8460 -26 8532 -17
rect 8460 -17 8532 -8
rect 8460 -8 8532 0
rect 8460 0 8532 8
rect 8460 8 8532 17
rect 8460 17 8532 26
rect 8460 26 8532 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 8316 316 8388 325
rect 8316 325 8388 334
rect 8316 334 8388 343
rect 8316 343 8388 352
rect 8316 352 8388 360
rect 8316 360 8388 369
rect 8316 369 8388 378
rect 8316 378 8388 387
rect 8388 316 8460 325
rect 8388 325 8460 334
rect 8388 334 8460 343
rect 8388 343 8460 352
rect 8388 352 8460 360
rect 8388 360 8460 369
rect 8388 369 8460 378
rect 8388 378 8460 387
rect 8460 316 8532 325
rect 8460 325 8532 334
rect 8460 334 8532 343
rect 8460 343 8532 352
rect 8460 352 8532 360
rect 8460 360 8532 369
rect 8460 369 8532 378
rect 8460 378 8532 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 8316 668 8388 677
rect 8316 677 8388 686
rect 8316 686 8388 695
rect 8316 695 8388 704
rect 8316 704 8388 712
rect 8316 712 8388 721
rect 8316 721 8388 730
rect 8316 730 8388 739
rect 8388 668 8460 677
rect 8388 677 8460 686
rect 8388 686 8460 695
rect 8388 695 8460 704
rect 8388 704 8460 712
rect 8388 712 8460 721
rect 8388 721 8460 730
rect 8388 730 8460 739
rect 8460 668 8532 677
rect 8460 677 8532 686
rect 8460 686 8532 695
rect 8460 695 8532 704
rect 8460 704 8532 712
rect 8460 712 8532 721
rect 8460 721 8532 730
rect 8460 730 8532 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< v2 >>
rect 8316 -35 8388 -26
rect 8316 -26 8388 -17
rect 8316 -17 8388 -8
rect 8316 -8 8388 0
rect 8316 0 8388 8
rect 8316 8 8388 17
rect 8316 17 8388 26
rect 8316 26 8388 35
rect 8388 -35 8460 -26
rect 8388 -26 8460 -17
rect 8388 -17 8460 -8
rect 8388 -8 8460 0
rect 8388 0 8460 8
rect 8388 8 8460 17
rect 8388 17 8460 26
rect 8388 26 8460 35
rect 8460 -35 8532 -26
rect 8460 -26 8532 -17
rect 8460 -17 8532 -8
rect 8460 -8 8532 0
rect 8460 0 8532 8
rect 8460 8 8532 17
rect 8460 17 8532 26
rect 8460 26 8532 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 8316 316 8388 325
rect 8316 325 8388 334
rect 8316 334 8388 343
rect 8316 343 8388 352
rect 8316 352 8388 360
rect 8316 360 8388 369
rect 8316 369 8388 378
rect 8316 378 8388 387
rect 8388 316 8460 325
rect 8388 325 8460 334
rect 8388 334 8460 343
rect 8388 343 8460 352
rect 8388 352 8460 360
rect 8388 360 8460 369
rect 8388 369 8460 378
rect 8388 378 8460 387
rect 8460 316 8532 325
rect 8460 325 8532 334
rect 8460 334 8532 343
rect 8460 343 8532 352
rect 8460 352 8532 360
rect 8460 360 8532 369
rect 8460 369 8532 378
rect 8460 378 8532 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 8316 668 8388 677
rect 8316 677 8388 686
rect 8316 686 8388 695
rect 8316 695 8388 704
rect 8316 704 8388 712
rect 8316 712 8388 721
rect 8316 721 8388 730
rect 8316 730 8388 739
rect 8388 668 8460 677
rect 8388 677 8460 686
rect 8388 686 8460 695
rect 8388 695 8460 704
rect 8388 704 8460 712
rect 8388 712 8460 721
rect 8388 721 8460 730
rect 8388 730 8460 739
rect 8460 668 8532 677
rect 8460 677 8532 686
rect 8460 686 8532 695
rect 8460 695 8532 704
rect 8460 704 8532 712
rect 8460 712 8532 721
rect 8460 721 8532 730
rect 8460 730 8532 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< viali >>
rect 8316 -35 8388 -26
rect 8316 -26 8388 -17
rect 8316 -17 8388 -8
rect 8316 -8 8388 0
rect 8316 0 8388 8
rect 8316 8 8388 17
rect 8316 17 8388 26
rect 8316 26 8388 35
rect 8388 -35 8460 -26
rect 8388 -26 8460 -17
rect 8388 -17 8460 -8
rect 8388 -8 8460 0
rect 8388 0 8460 8
rect 8388 8 8460 17
rect 8388 17 8460 26
rect 8388 26 8460 35
rect 8460 -35 8532 -26
rect 8460 -26 8532 -17
rect 8460 -17 8532 -8
rect 8460 -8 8532 0
rect 8460 0 8532 8
rect 8460 8 8532 17
rect 8460 17 8532 26
rect 8460 26 8532 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 8316 316 8388 325
rect 8316 325 8388 334
rect 8316 334 8388 343
rect 8316 343 8388 352
rect 8316 352 8388 360
rect 8316 360 8388 369
rect 8316 369 8388 378
rect 8316 378 8388 387
rect 8388 316 8460 325
rect 8388 325 8460 334
rect 8388 334 8460 343
rect 8388 343 8460 352
rect 8388 352 8460 360
rect 8388 360 8460 369
rect 8388 369 8460 378
rect 8388 378 8460 387
rect 8460 316 8532 325
rect 8460 325 8532 334
rect 8460 334 8532 343
rect 8460 343 8532 352
rect 8460 352 8532 360
rect 8460 360 8532 369
rect 8460 369 8532 378
rect 8460 378 8532 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 8316 668 8388 677
rect 8316 677 8388 686
rect 8316 686 8388 695
rect 8316 695 8388 704
rect 8316 704 8388 712
rect 8316 712 8388 721
rect 8316 721 8388 730
rect 8316 730 8388 739
rect 8388 668 8460 677
rect 8388 677 8460 686
rect 8388 686 8460 695
rect 8388 695 8460 704
rect 8388 704 8460 712
rect 8388 712 8460 721
rect 8388 721 8460 730
rect 8388 730 8460 739
rect 8460 668 8532 677
rect 8460 677 8532 686
rect 8460 686 8532 695
rect 8460 695 8532 704
rect 8460 704 8532 712
rect 8460 712 8532 721
rect 8460 721 8532 730
rect 8460 730 8532 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< m3 >>
rect 108 -44 8676 44
rect 108 -44 8676 44
rect 8604 44 8676 132
rect 108 132 8316 220
rect 8388 132 8532 220
rect 8604 132 8676 220
rect 108 220 180 308
rect 8604 220 8676 308
rect 108 308 180 396
rect 252 308 324 396
rect 396 308 8676 396
rect 108 396 180 484
rect 8604 396 8676 484
rect 108 484 8532 572
rect 8604 484 8676 572
rect 108 572 180 660
rect 8604 572 8676 660
rect 108 660 180 748
rect 252 660 8676 748
rect 108 748 180 836
rect 108 836 8676 924
rect 108 836 8676 924
<< rm3 >>
rect 8316 132 8388 220
rect 324 308 396 396
<< labels >>
flabel m3 s 108 -44 8676 44 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 108 836 8676 924 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 8712 0 1056
<< end >>
