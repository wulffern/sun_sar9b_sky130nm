
*-------------------------------------------------------------
* SUNSAR_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNSAR_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNSAR_NCHDLR <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_NCHDLR D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNSAR_RM1 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_RM1 A B
R1 A B 1m
.ENDS

*-------------------------------------------------------------
* SUNSAR_CAP_BSSW_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_CAP_BSSW_CV A B
C1 A B 100f
.ENDS

*-------------------------------------------------------------
* SUNSAR_CAP_BSSW5_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_CAP_BSSW5_CV A B
XCAPB0 A B SUNSAR_CAP_BSSW_CV
XCAPB1 A B SUNSAR_CAP_BSSW_CV
XCAPB2 A B SUNSAR_CAP_BSSW_CV
XCAPB3 A B SUNSAR_CAP_BSSW_CV
XCAPB4 A B SUNSAR_CAP_BSSW_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_TIEH_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_TIEH_CV Y BULKP BULKN AVDD AVSS
XMN0 A A AVSS BULKN SUNSAR_NCHDL
XMP0 Y A AVDD BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_TIEL_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_TIEL_CV Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNSAR_NCHDL
XMP0 A A AVDD BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_TAPCELLB_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNSAR_NCHDL
XMP1 AVDD AVDD AVDD AVDD SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_IVX1_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNSAR_NCHDL
XMP0 Y A AVDD BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_IVX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_IVX4_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNSAR_NCHDL
XMN1 AVSS A Y BULKN SUNSAR_NCHDL
XMN2 Y A AVSS BULKN SUNSAR_NCHDL
XMN3 AVSS A Y BULKN SUNSAR_NCHDL
XMP0 Y A AVDD BULKP SUNSAR_PCHDL
XMP1 AVDD A Y BULKP SUNSAR_PCHDL
XMP2 Y A AVDD BULKP SUNSAR_PCHDL
XMP3 AVDD A Y BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_BFX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_BFX1_CV A Y BULKP BULKN AVDD AVSS
XMN0 AVSS A B BULKN SUNSAR_NCHDL
XMN1 Y B AVSS BULKN SUNSAR_NCHDL
XMP0 AVDD A B BULKP SUNSAR_PCHDL
XMP1 Y B AVDD BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_NRX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_NRX1_CV A B Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNSAR_NCHDL
XMN1 AVSS B Y BULKN SUNSAR_NCHDL
XMP0 N1 A AVDD BULKP SUNSAR_PCHDL
XMP1 Y B N1 BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_NDX1_CV A B Y BULKP BULKN AVDD AVSS
XMN0 N1 A AVSS BULKN SUNSAR_NCHDL
XMN1 Y B N1 BULKN SUNSAR_NCHDL
XMP0 Y A AVDD BULKP SUNSAR_PCHDL
XMP1 AVDD B Y BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_ORX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_ORX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNSAR_NRX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNSAR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_ANX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_ANX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNSAR_NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNSAR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_IVTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_IVTRIX1_CV A C CN Y BULKP BULKN AVDD AVSS
XMN0 N1 A AVSS BULKN SUNSAR_NCHDL
XMN1 Y C N1 BULKN SUNSAR_NCHDL
XMP0 N2 A AVDD BULKP SUNSAR_PCHDL
XMP1 Y CN N2 BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_NDTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_NDTRIX1_CV A C CN RN Y BULKP BULKN AVDD AVSS
XMN2 N1 RN AVSS BULKN SUNSAR_NCHDL
XMN0 N2 A N1 BULKN SUNSAR_NCHDL
XMN1 Y C N2 BULKN SUNSAR_NCHDL
XMP2 AVDD RN N2 BULKP SUNSAR_PCHDL
XMP0 N2 A AVDD BULKP SUNSAR_PCHDL
XMP1 Y CN N2 BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_DFRNQNX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS SUNSAR_TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS AVDD AVSS SUNSAR_NDX1_CV
XA2 CKN CKB AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS AVDD AVSS SUNSAR_IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS AVDD AVSS SUNSAR_IVTRIX1_CV
XA5 A0 A1 AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS AVDD AVSS SUNSAR_IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS AVDD AVSS SUNSAR_NDTRIX1_CV
XA8 QN Q AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_SWX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SWX4_CV A Y VREF AVSS BULKP BULKN
XMN0 Y A AVSS BULKN SUNSAR_NCHDL
XMN1 AVSS A Y BULKN SUNSAR_NCHDL
XMN2 Y A AVSS BULKN SUNSAR_NCHDL
XMN3 AVSS A Y BULKN SUNSAR_NCHDL
XMP0 Y A VREF BULKP SUNSAR_PCHDL
XMP1 VREF A Y BULKP SUNSAR_PCHDL
XMP2 Y A VREF BULKP SUNSAR_PCHDL
XMP3 VREF A Y BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_TGPD_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_TGPD_CV C A B BULKP BULKN AVDD AVSS
XMN0 AVSS C CN BULKN SUNSAR_NCHDL
XMN1 B C AVSS BULKN SUNSAR_NCHDL
XMN2 A CN B BULKN SUNSAR_NCHDL
XMP0 AVDD C CN BULKP SUNSAR_PCHDL
XMP1_DMY B AVDD AVDD BULKP SUNSAR_PCHDL
XMP2 A C B BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_SAREMX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SAREMX1_CV A B EN ENO RST_N BULKP BULKN AVDD AVSS
XMN0 N3 EN AM BULKN SUNSAR_NCHDL
XMN1 N3 B AVSS BULKN SUNSAR_NCHDL
XMN2 AVSS A N3 BULKN SUNSAR_NCHDL
XMN3 ENO AM AVSS BULKN SUNSAR_NCHDL
XMP0 AVDD RST_N AM BULKP SUNSAR_PCHDL
XMP1 N2 B ENO BULKP SUNSAR_PCHDL
XMP2 N1 A N2 BULKP SUNSAR_PCHDL
XMP3 AVDD AM N1 BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARLTX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARLTX1_CV A CHL RST_N EN LCK_N BULKP BULKN AVDD AVSS
XMN0 N1 A AVSS BULKN SUNSAR_NCHDL
XMN1 N3 LCK_N N1 BULKN SUNSAR_NCHDL
XMN2 CHL EN N3 BULKN SUNSAR_NCHDL
XMP0 NP2 RST_N AVDD BULKP SUNSAR_PCHDL
XMP1 NP1 RST_N NP2 BULKP SUNSAR_PCHDL
XMP2 CHL RST_N NP1 BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARCEX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARCEX1_CV A B Y RST BULKP BULKN AVDD AVSS
XMN0 N4 RST AVSS BULKN SUNSAR_NCHDL
XMN1 AVSS RST N4 BULKN SUNSAR_NCHDL
XMN2 N1 RST AVSS BULKN SUNSAR_NCHDL
XMN3 Y RST N1 BULKN SUNSAR_NCHDL
XMP0 N2 A Y BULKP SUNSAR_PCHDL
XMP1 AVDD A N2 BULKP SUNSAR_PCHDL
XMP2 N3 B AVDD BULKP SUNSAR_PCHDL
XMP3 Y B N3 BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARCMPHX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARCMPHX1_CV CI CK CO VMR N1 N2 BULKP BULKN AVDD AVSS
XMN0 N1 CK AVSS BULKN SUNSAR_NCHDL
XMN1 N2 CI N1 BULKN SUNSAR_NCHDL
XMN2 N1 CI N2 BULKN SUNSAR_NCHDL
XMN3 N2 CI N1 BULKN SUNSAR_NCHDL
XMN4 N1 CI N2 BULKN SUNSAR_NCHDL
XMN5 N2 CI N1 BULKN SUNSAR_NCHDL
XMN6 CO VMR N2 BULKN SUNSAR_NCHDL
XMP0 AVDD CK N1 BULKP SUNSAR_PCHDL
XMP1 N2 CK AVDD BULKP SUNSAR_PCHDL
XMP2 AVDD AVDD N2 BULKP SUNSAR_PCHDL
XMP3 CO CK AVDD BULKP SUNSAR_PCHDL
XMP4 AVDD VMR CO BULKP SUNSAR_PCHDL
XMP5 CO VMR AVDD BULKP SUNSAR_PCHDL
XMP6 AVDD VMR CO BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARKICKHX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARKICKHX1_CV CI CK CKN BULKP BULKN AVDD AVSS
XMN0 N1 CKN AVSS BULKN SUNSAR_NCHDL
XMN1 N1 CI N1 BULKN SUNSAR_NCHDL
XMN2 N1 CI N1 BULKN SUNSAR_NCHDL
XMN3 N1 CI N1 BULKN SUNSAR_NCHDL
XMN4 N1 CI N1 BULKN SUNSAR_NCHDL
XMN5 N1 CI N1 BULKN SUNSAR_NCHDL
XMN6 AVDD CK N1 BULKN SUNSAR_NCHDL
XMP0 AVDD CKN N1 BULKP SUNSAR_PCHDL
XMP1_DMY AVDD AVDD AVDD BULKP SUNSAR_PCHDL
XMP2_DMY AVDD AVDD AVDD BULKP SUNSAR_PCHDL
XMP3_DMY AVDD AVDD AVDD BULKP SUNSAR_PCHDL
XMP4_DMY AVDD AVDD AVDD BULKP SUNSAR_PCHDL
XMP5_DMY AVDD AVDD AVDD BULKP SUNSAR_PCHDL
XMP6_DMY AVDD AVDD AVDD BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARBSSWCTRL_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARBSSWCTRL_CV C GN GNG TIE_H BULKP BULKN AVDD AVSS
XMN0 N1 C AVSS BULKN SUNSAR_NCHDL
XMN1 GN TIE_H N1 BULKN SUNSAR_NCHDL
XMP0 GNG C GN BULKP SUNSAR_PCHDL
XMP1 AVDD GN GNG BULKP SUNSAR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_CAP32C_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_CAP32C_CV C1A C1B C2 C4 C8 C16 CTOP AVSS
C1 C1A CTOP 0.2f
C2 C1B CTOP 0.2f
C3 C2 CTOP 0.4f
C4 C4 CTOP 0.8f
C5 C8 CTOP 1.6f
C6 C16 CTOP 3.2f
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARCMPX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARCMPX1_CV CPI CNI CPO CNO CK_CMP CK_SAMPLE DONE AVDD AVSS
XA0 AVDD AVSS SUNSAR_TAPCELLB_CV
XA1 CPI CK_B CK_N AVDD AVSS AVDD AVSS SUNSAR_SARKICKHX1_CV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS AVDD AVSS SUNSAR_SARCMPHX1_CV
XA2a CPO_I CPO AVDD AVSS AVDD AVSS SUNSAR_IVX4_CV
XA3a CNO_I CNO AVDD AVSS AVDD AVSS SUNSAR_IVX4_CV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS AVDD AVSS SUNSAR_SARCMPHX1_CV
XA4 CNI CK_B CK_N AVDD AVSS AVDD AVSS SUNSAR_SARKICKHX1_CV
XA9 CK_N CK_B AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA10 DONE_N CK_A CK_N AVDD AVSS AVDD AVSS SUNSAR_NDX1_CV
XA11 CK_SAMPLE DONE DONE_N AVDD AVSS AVDD AVSS SUNSAR_NRX1_CV
XA12 CK_CMP CK_A AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA13 AVDD AVSS SUNSAR_TAPCELLB_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARBSSW_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARBSSW_CV VI CK CKN TIE_L VO1 VO2 AVDD AVSS
XM1 VI GN VO1 AVSS SUNSAR_NCHDLR
XM2 VI GN VO1 AVSS SUNSAR_NCHDLR
XM3 VI GN VO1 AVSS SUNSAR_NCHDLR
XM4 VI GN VO1 AVSS SUNSAR_NCHDLR
XM5 VI TIE_L VO2 AVSS SUNSAR_NCHDLR
XM6 VI TIE_L VO2 AVSS SUNSAR_NCHDLR
XM7 VI TIE_L VO2 AVSS SUNSAR_NCHDLR
XM8 VI TIE_L VO2 AVSS SUNSAR_NCHDLR
XA5b AVDD AVSS SUNSAR_TAPCELLB_CV
XA0 CK CKN AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA3 CKN VI VS AVDD AVSS AVDD AVSS SUNSAR_TGPD_CV
XA4 CKN GN GNG TIE_H AVDD AVSS AVDD AVSS SUNSAR_SARBSSWCTRL_CV
XA1 TIE_H AVDD AVSS AVDD AVSS SUNSAR_TIEH_CV
XA7 AVDD AVSS SUNSAR_TAPCELLB_CV
XA2 TIE_L AVDD AVSS AVDD AVSS SUNSAR_TIEL_CV
XA5 AVDD AVSS SUNSAR_TAPCELLB_CV
XCAPB1 GNG VS SUNSAR_CAP_BSSW5_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARMRYX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARMRYX1_CV CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS
XA0 AVDD AVSS SUNSAR_TAPCELLB_CV
XA1 CMP_OP CMP_ON EN ENO RST_N AVDD AVSS AVDD AVSS SUNSAR_SAREMX1_CV
XA2 ENO LCK_N AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA4 CMP_OP CHL_OP RST_N EN LCK_N AVDD AVSS AVDD AVSS SUNSAR_SARLTX1_CV
XA5 CMP_ON CHL_ON RST_N EN LCK_N AVDD AVSS AVDD AVSS SUNSAR_SARLTX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARDIGEX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARDIGEX4_CV CMP_OP CMP_ON EN RST_N ENO DONE CP0 CP1 CN0 CN1 CEIN CEO CKS VREF AVDD AVSS
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS SUNSAR_SARMRYX1_CV
XA2 CHL_ON CN1 VREF AVSS AVDD AVSS SUNSAR_SWX4_CV
XA3 CN1 CP1 VREF AVSS AVDD AVSS SUNSAR_SWX4_CV
XA4 CHL_OP CP0 VREF AVSS AVDD AVSS SUNSAR_SWX4_CV
XA5 CP0 CN0 VREF AVSS AVDD AVSS SUNSAR_SWX4_CV
XA6 CN0 CP1 CE CKS AVDD AVSS AVDD AVSS SUNSAR_SARCEX1_CV
XA7 ENO ENO_N AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA8 ENO_N DONE AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA9 ENO_N CE CE1 AVDD AVSS AVDD AVSS SUNSAR_NDX1_CV
XA10 CE1 CE1_N AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA11 CE1_N CEIN CEO1 AVDD AVSS AVDD AVSS SUNSAR_NRX1_CV
XA12 CEO1 CEO AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA13 AVDD AVSS SUNSAR_TAPCELLB_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_CDAC8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_CDAC8_CV CP_11 CP_10 CP_9 CP_8 CP_7 CP_6 CP_5 CP_4 CP_3 CP_2 CP_1 CP_0 CTOP AVSS
XC1 CP_10 CP_10 CP_10 CP_10 CP_10 CP_10 CTOP AVSS SUNSAR_CAP32C_CV
XC64a<0> CP_8 CP_8 CP_8 CP_8 CP_8 CP_8 CTOP AVSS SUNSAR_CAP32C_CV
XC32a<0> AVSS CP_0 CP_1 CP_2 CP_3 CP_7 CTOP AVSS SUNSAR_CAP32C_CV
XC128a<1> CP_11 CP_11 CP_11 CP_11 CP_11 CP_11 CTOP AVSS SUNSAR_CAP32C_CV
XC128b<2> CP_10 CP_10 CP_10 CP_10 CP_10 CP_10 CTOP AVSS SUNSAR_CAP32C_CV
X16ab CP_5 CP_5 CP_5 CP_5 CP_4 CP_6 CTOP AVSS SUNSAR_CAP32C_CV
XC64b<1> CP_9 CP_9 CP_9 CP_9 CP_9 CP_9 CTOP AVSS SUNSAR_CAP32C_CV
XC0 CP_11 CP_11 CP_11 CP_11 CP_11 CP_11 CTOP AVSS SUNSAR_CAP32C_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_CDAC7_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_CDAC7_CV CP_9 CP_8 CP_7 CP_6 CP_5 CP_4 CP_3 CP_2 CP_1 CP_0 CTOP AVSS
XC1 CP_8 CP_8 CP_8 CP_8 CP_8 CP_8 CTOP AVSS SUNSAR_CAP32C_CV
XC32a<0> AVSS CP_0 CP_1 CP_2 CP_3 CP_7 CTOP AVSS SUNSAR_CAP32C_CV
X16ab CP_5 CP_5 CP_5 CP_5 CP_4 CP_6 CTOP AVSS SUNSAR_CAP32C_CV
XC0 CP_9 CP_9 CP_9 CP_9 CP_9 CP_9 CTOP AVSS SUNSAR_CAP32C_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_SAR9B_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D_8 D_7 D_6 D_5 D_4 D_3 D_2 D_1 D_0 EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
XB1 SAR_IP CK_SAMPLE_BSSW NCCA CEIN SARP SARN AVDD AVSS SUNSAR_SARBSSW_CV
XB2 SAR_IN CK_SAMPLE_BSSW NCCB CEIN SARN SARP AVDD AVSS SUNSAR_SARBSSW_CV
XDAC1 CP_11 CP_10 D_7 CP_8 D_6 CP_6 D_5 CP_4 D_4 D_3 D_2 D_1 SARP AVSS SUNSAR_CDAC8_CV
XDAC2 D_8 CN_10 CN_9 CN_8 CN_7 CN_6 CN_5 CN_4 CN_3 CN_2 CN_1 CN_0 SARN AVSS SUNSAR_CDAC8_CV
XA0 CMP_OP CMP_ON EN EN ENO0 DONE0 CP_10 CP_11 CN_10 D_8 CEIN CEO0 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA1 CMP_OP CMP_ON ENO0 EN ENO1 DONE1 CP_8 D_7 CN_8 CN_9 CEO0 CEO1 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA2 CMP_OP CMP_ON ENO1 EN ENO2 DONE2 CP_6 D_6 CN_6 CN_7 CEO1 CEO2 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA3 CMP_OP CMP_ON ENO2 EN ENO3 DONE3 CP_4 D_5 CN_4 CN_5 CEO2 CEO3 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA4 CMP_OP CMP_ON ENO3 EN ENO4 DONE4 NC2A D_4 CN_3 NC2B CEO3 CEO4 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA5 CMP_OP CMP_ON ENO4 EN ENO5 DONE5 NC3A D_3 CN_2 NC3B CEO4 CEO5 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA6 CMP_OP CMP_ON ENO5 EN ENO6 DONE6 NC4A D_2 CN_1 NC4B CEO5 CEO6 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA7 CMP_OP CMP_ON ENO6 EN ENO7 DONE7 NC5A D_1 CN_0 NC5B CEO6 CEO7 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA8 CMP_OP CMP_ON ENO7 EN ENO8 DONE NC6A D_0 NC6C NC6B CEO7 CK_CMP CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA20 SARP SARN CMP_OP CMP_ON CK_CMP CK_SAMPLE DONE AVDD AVSS SUNSAR_SARCMPX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_SAR8B_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SAR8B_CV SAR_IP SAR_IN SARN SARP DONE D_7 D_6 D_5 D_4 D_3 D_2 D_1 D_0 EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
XB1 SAR_IP CK_SAMPLE_BSSW NCCA CEIN SARP SARN AVDD AVSS SUNSAR_SARBSSW_CV
XB2 SAR_IN CK_SAMPLE_BSSW NCCB CEIN SARN SARP AVDD AVSS SUNSAR_SARBSSW_CV
XDAC1 CP_9 CP_8 D_6 CP_6 D_5 CP_4 D_4 D_3 D_2 D_1 SARP AVSS SUNSAR_CDAC7_CV
XDAC2 D_7 CN_8 CN_7 CN_6 CN_5 CN_4 CN_3 CN_2 CN_1 CN_0 SARN AVSS SUNSAR_CDAC7_CV
XA0 CMP_OP CMP_ON EN EN ENO0 DONE0 CP_8 CP_9 CN_8 D_7 CEIN CEO0 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA1 CMP_OP CMP_ON ENO0 EN ENO1 DONE1 CP_6 D_6 CN_6 CN_7 CEO0 CEO1 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA2 CMP_OP CMP_ON ENO1 EN ENO2 DONE2 CP_4 D_5 CN_4 CN_5 CEO1 CEO2 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA3 CMP_OP CMP_ON ENO2 EN ENO3 DONE3 NC2A D_4 CN_3 NC2B CEO2 CEO3 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA4 CMP_OP CMP_ON ENO3 EN ENO4 DONE4 NC3A D_3 CN_2 NC3B CEO3 CEO4 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA5 CMP_OP CMP_ON ENO4 EN ENO5 DONE5 NC4A D_2 CN_1 NC4B CEO4 CEO5 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA6 CMP_OP CMP_ON ENO5 EN ENO6 DONE6 NC5A D_1 CN_0 NC5B CEO5 CEO6 CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA7 CMP_OP CMP_ON ENO6 EN ENO7 DONE NC6A D_0 NC6C NC6B CEO6 CK_CMP CK_SAMPLE VREF AVDD AVSS SUNSAR_SARDIGEX4_CV
XA20 SARP SARN CMP_OP CMP_ON CK_CMP CK_SAMPLE DONE AVDD AVSS SUNSAR_SARCMPX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_SARCAPTURE_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_SARCAPTURE_CV CKS ENABLE CK_SAMPLE CK_SAMPLE_BSSW EN D_7 D_6 D_5 D_4 D_3 D_2 D_1 D_0 DO_7 DO_6 DO_5 DO_4 DO_3 DO_2 DO_1 DO_0 DONE AVDD AVSS
XB07 D_7 DONE ENABLE_B DO_7 DN7 AVDD AVSS SUNSAR_DFRNQNX1_CV
XC08 D_6 DONE ENABLE_B DO_6 DN6 AVDD AVSS SUNSAR_DFRNQNX1_CV
XD09 D_5 DONE ENABLE_B DO_5 DN5 AVDD AVSS SUNSAR_DFRNQNX1_CV
XE10 D_4 DONE ENABLE_B DO_4 DN4 AVDD AVSS SUNSAR_DFRNQNX1_CV
XF11 D_3 DONE ENABLE_B DO_3 DN3 AVDD AVSS SUNSAR_DFRNQNX1_CV
XG12 D_2 DONE ENABLE_B DO_2 DN2 AVDD AVSS SUNSAR_DFRNQNX1_CV
XH13 D_1 DONE ENABLE_B DO_1 DN1 AVDD AVSS SUNSAR_DFRNQNX1_CV
XI14 D_0 DONE ENABLE_B DO_0 DM0 AVDD AVSS SUNSAR_DFRNQNX1_CV
XA1 AVDD AVSS SUNSAR_TAPCELLB_CV
XA2 ENABLE ENABLE_N AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA3 ENABLE_N ENABLE_B AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA4 CKS CKS_B AVDD AVSS AVDD AVSS SUNSAR_BFX1_CV
XA5 CKS_B ENABLE_N CK_SAMPLE AVDD AVSS AVDD AVSS SUNSAR_ORX1_CV
XA5a CK_SAMPLE EN AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA6 CKS_B ENABLE_B CK_SAMPLE_BSSW AVDD AVSS AVDD AVSS SUNSAR_ANX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_DFQNX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_DFQNX1_CV D CK Q QN AVDD AVSS
XA0 AVDD AVSS SUNSAR_TAPCELLB_CV
XA1 CK CKN AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA2 CKN CKB AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS AVDD AVSS SUNSAR_IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS AVDD AVSS SUNSAR_IVTRIX1_CV
XA5 A0 A1 AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS AVDD AVSS SUNSAR_IVTRIX1_CV
XA7 Q CKN CKB QN AVDD AVSS AVDD AVSS SUNSAR_IVTRIX1_CV
XA8 QN Q AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNSAR_CAPT8B_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_CAPT8B_CV CKS ENABLE CK_SAMPLE CK_SAMPLE_BSSW EN D_7 D_6 D_5 D_4 D_3 D_2 D_1 D_0 DO_7 DO_6 DO_5 DO_4 DO_3 DO_2 DO_1 DO_0 DONE AVDD AVSS TIE_L
XB07 D_7 DONE DO_7 DN7 AVDD AVSS SUNSAR_DFQNX1_CV
XC08 D_6 DONE DO_6 DN6 AVDD AVSS SUNSAR_DFQNX1_CV
XD09 D_5 DONE DO_5 DN5 AVDD AVSS SUNSAR_DFQNX1_CV
XE10 D_4 DONE DO_4 DN4 AVDD AVSS SUNSAR_DFQNX1_CV
XF11 D_3 DONE DO_3 DN3 AVDD AVSS SUNSAR_DFQNX1_CV
XG12 D_2 DONE DO_2 DN2 AVDD AVSS SUNSAR_DFQNX1_CV
XH13 D_1 DONE DO_1 DN1 AVDD AVSS SUNSAR_DFQNX1_CV
XI14 D_0 DONE DO_0 DM0 AVDD AVSS SUNSAR_DFQNX1_CV
XA1 AVDD AVSS SUNSAR_TAPCELLB_CV
XA2 ENABLE ENABLE_N AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA3 ENABLE_N ENABLE_B AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA4 CKS CKS_B AVDD AVSS AVDD AVSS SUNSAR_BFX1_CV
XA5 CKS_B ENABLE_N CK_SAMPLE AVDD AVSS AVDD AVSS SUNSAR_ORX1_CV
XA5a CK_SAMPLE EN AVDD AVSS AVDD AVSS SUNSAR_IVX1_CV
XA6 CKS_B ENABLE_B CK_SAMPLE_BSSW AVDD AVSS AVDD AVSS SUNSAR_ANX1_CV
XA2 TIE_L AVDD AVSS AVDD AVSS SUNSAR_TIEL_CV
.ENDS
