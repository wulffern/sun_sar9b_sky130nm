magic
tech sky130A
timestamp 1712959200
<< checkpaint >>
rect 0 0 1260 440
<< locali >>
rect 378 379 828 413
rect 199 193 233 369
rect 415 291 449 325
rect 415 203 449 237
rect 162 159 270 193
rect -54 66 54 110
rect 199 71 233 159
rect 415 115 449 149
rect 516 61 550 379
rect 811 291 845 325
rect 1027 281 1061 369
rect 990 247 1098 281
rect 811 203 845 237
rect 811 115 845 149
rect 1027 105 1061 193
rect 990 71 1098 105
rect 1206 66 1314 110
rect 516 27 828 61
<< metal3 >>
rect 378 0 470 440
rect 774 0 866 440
use SUNSAR_NCHDL  MN0
timestamp 1712959200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_NCHDL  MN1
timestamp 1712959200
transform 1 0 0 0 1 88
box -90 -66 630 242
use SUNSAR_NCHDL  MN2
timestamp 1712959200
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNSAR_NCHDL  MN3
timestamp 1712959200
transform 1 0 0 0 1 264
box -90 -66 630 242
use SUNSAR_PCHDL  MP0
timestamp 1712959200
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_PCHDL  MP1
timestamp 1712959200
transform 1 0 630 0 1 88
box 0 -66 720 242
use SUNSAR_PCHDL  MP2
timestamp 1712959200
transform 1 0 630 0 1 176
box 0 -66 720 242
use SUNSAR_PCHDL  MP3
timestamp 1712959200
transform 1 0 630 0 1 264
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1712959200
transform 1 0 774 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1712959200
transform 1 0 774 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut2
timestamp 1712959200
transform 1 0 378 0 1 27
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut3
timestamp 1712959200
transform 1 0 378 0 1 203
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut4
timestamp 1712959200
transform 1 0 378 0 1 203
box 0 0 92 34
<< labels >>
flabel locali s 990 71 1098 105 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 990 247 1098 281 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 162 159 270 193 0 FreeSans 400 0 0 0 RST
port 4 nsew signal bidirectional
flabel locali s 378 379 486 413 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 5 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 6 nsew signal bidirectional
flabel metal3 s 774 0 866 440 0 FreeSans 400 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel metal3 s 378 0 470 440 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 440
<< end >>
