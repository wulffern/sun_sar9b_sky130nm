magic
tech sky130A
magscale 1 2
timestamp 1712087342
<< locali >>
rect 19026 32668 19242 32736
rect 162 31524 378 31592
rect 1818 27476 2034 27544
rect 10206 2518 10422 2586
rect 10206 1110 10422 1178
<< metal1 >>
rect -1922 -1796 -1854 37062
rect -1710 36878 24066 37062
rect -1710 36158 24066 36342
rect -1710 -1256 -1526 36158
rect -990 35438 23346 35622
rect -990 15254 -806 35438
rect 3114 34428 3518 34496
rect 8154 34428 8558 34496
rect 13194 34428 13598 34496
rect 3450 33928 3518 34428
rect 5134 33928 5202 34056
rect 3450 33860 5202 33928
rect 8490 33928 8558 34428
rect 10174 33928 10242 34056
rect 8490 33860 10242 33928
rect 13530 33928 13598 34428
rect 15214 33928 15282 34056
rect 13530 33860 15282 33928
rect 9132 18586 9200 20446
rect 9320 18586 9388 21748
rect 9508 18586 9576 20632
rect 9696 18586 9764 21934
rect 9884 18586 9952 20818
rect 10072 18586 10140 22120
rect 10260 18586 10328 21004
rect 10448 18586 10516 21190
rect 10636 18586 10704 21376
rect 10824 18586 10892 21562
rect 11464 18586 11532 23422
rect 11652 18586 11720 23236
rect 11840 18586 11908 23050
rect 12028 18586 12096 22864
rect 12216 18586 12284 22678
rect 12404 18586 12472 20260
rect 12592 18586 12660 22492
rect 12780 18586 12848 20074
rect 12968 18586 13036 22306
rect 13156 18586 13224 19888
rect 23162 15254 23346 35438
rect -990 15186 68 15254
rect 22288 15186 23346 15254
rect -990 11854 -806 15186
rect 23162 11854 23346 15186
rect -990 11786 68 11854
rect 22288 11786 23346 11854
rect -990 8454 -806 11786
rect 23162 8454 23346 11786
rect -990 8386 68 8454
rect 22288 8386 23346 8454
rect -990 5054 -806 8386
rect 23162 5054 23346 8386
rect -990 4986 68 5054
rect 22288 4986 23346 5054
rect -990 -536 -806 4986
rect 23162 -536 23346 4986
rect -990 -720 23346 -536
rect 23882 -1256 24066 36158
rect -1710 -1440 24066 -1256
rect 24210 -1584 24278 37062
rect -1710 -1652 24278 -1584
rect -1922 -1864 24278 -1796
<< metal2 >>
rect 1386 34462 1790 34530
rect 6426 34462 6830 34530
rect 11466 34462 11870 34530
rect 16506 34462 16910 34530
rect -1854 33988 162 34056
rect 1722 33928 1790 34462
rect 4270 33928 4338 34056
rect 1722 33860 4338 33928
rect 6762 33928 6830 34462
rect 9310 33928 9378 34056
rect 6762 33860 9378 33928
rect 11802 33928 11870 34462
rect 14350 33928 14418 34056
rect 11802 33860 14418 33928
rect 16842 33928 16910 34462
rect 18342 34428 19934 34496
rect 19390 33928 19458 34056
rect 16842 33860 19458 33928
rect 19866 33562 19934 34428
rect 19866 33494 20430 33562
rect 19302 33108 20430 33176
rect 19302 32736 19370 33108
rect 22086 32932 22322 33000
rect 702 32668 938 32736
rect 4014 32668 4250 32736
rect 5742 32668 5978 32736
rect 9054 32668 9290 32736
rect 10782 32668 11018 32736
rect 14094 32668 14330 32736
rect 15822 32668 16058 32736
rect 19134 32668 19370 32736
rect 19566 31876 19674 31944
rect 22254 31876 22322 32932
rect 19614 31808 22322 31876
rect 94 31464 162 31592
rect 4270 31464 4338 31592
rect 5134 31464 5202 31592
rect 9310 31464 9378 31592
rect 10174 31464 10242 31592
rect 14350 31464 14418 31592
rect 15214 31464 15282 31592
rect 19390 31464 19458 31592
rect 94 31396 19674 31464
rect 19734 28512 21606 28580
rect 162 27476 18018 27544
rect 19734 27192 19802 28512
rect 21546 28444 21654 28512
rect 94 26916 162 27192
rect 4270 26916 4338 27192
rect 5134 26916 5202 27192
rect 9310 26916 9378 27192
rect 10174 26916 10242 27192
rect 14350 26916 14418 27192
rect 15214 26916 15282 27192
rect 19390 26916 19458 27192
rect 19566 27124 19802 27192
rect 20206 27598 20862 27666
rect 94 26848 19674 26916
rect 126 26696 19642 26764
rect 126 26420 194 26696
rect 4270 26420 4338 26696
rect 5166 26420 5234 26696
rect 9310 26420 9378 26696
rect 10206 26420 10274 26696
rect 14350 26420 14418 26696
rect 15246 26420 15314 26696
rect 19390 26420 19458 26696
rect 20206 26556 20274 27598
rect 19582 26488 20274 26556
rect 19550 26420 19642 26488
rect 3418 25052 5234 25120
rect 3418 24992 3486 25052
rect 1418 24924 1790 24992
rect 3114 24924 3486 24992
rect 1722 24600 1790 24924
rect 4270 24600 4338 24728
rect 5166 24660 5234 25052
rect 8458 25052 10274 25120
rect 8458 24992 8526 25052
rect 6458 24924 6830 24992
rect 8154 24924 8526 24992
rect 1722 24532 4338 24600
rect 6762 24600 6830 24924
rect 9310 24600 9378 24728
rect 10206 24660 10274 25052
rect 13498 25052 15314 25120
rect 13498 24992 13566 25052
rect 11498 24924 11870 24992
rect 13194 24924 13566 24992
rect 6762 24532 9378 24600
rect 11802 24600 11870 24924
rect 14350 24600 14418 24728
rect 15246 24660 15314 25052
rect 18538 24992 18606 25052
rect 16538 24924 16910 24992
rect 18234 24924 18606 24992
rect 11802 24532 14418 24600
rect 16842 24600 16910 24924
rect 19390 24600 19458 24728
rect 16842 24532 19458 24600
rect 11464 23422 16372 23490
rect 11652 23236 13612 23304
rect 11264 23050 11908 23118
rect 8504 22864 12096 22932
rect 6224 22678 12284 22746
rect 3464 22492 12660 22560
rect 1184 22306 13036 22374
rect 6067 22120 10140 22188
rect 3620 21934 9764 22002
rect 1027 21748 9388 21816
rect 10824 21562 16072 21630
rect 10636 21376 13911 21444
rect 10448 21190 11032 21258
rect 8803 21004 10328 21072
rect 5924 20818 9952 20886
rect 3763 20632 9576 20700
rect 884 20446 9200 20514
rect 5234 20260 12472 20328
rect 4338 20074 12848 20142
rect 194 19888 13224 19956
rect 8580 18654 8648 19584
rect 20322 19516 20390 19856
rect 13708 18654 13776 19212
rect 20598 19144 20666 19856
rect 10314 2518 10550 2586
rect 10482 1178 10550 2518
rect 10482 1110 12042 1178
rect 9272 -1652 9340 562
rect 13016 -1652 13084 562
<< metal3 >>
rect 194 19956 262 28708
rect 594 24166 778 35622
rect 884 20514 952 28738
rect 1027 21816 1095 29618
rect 1184 22374 1252 30498
rect 1386 24166 1570 36342
rect 1962 28092 2146 37062
rect 2570 28092 2754 37062
rect 3146 24166 3330 36342
rect 3464 22560 3532 30498
rect 3620 22002 3688 29618
rect 3763 20700 3831 28738
rect 3938 24166 4122 35622
rect 4338 20142 4406 28708
rect 5234 20328 5302 28708
rect 5634 24166 5818 35622
rect 5924 20886 5992 28738
rect 6067 22188 6135 29618
rect 6224 22746 6292 30498
rect 6426 24166 6610 36342
rect 7002 28092 7186 37062
rect 7610 28092 7794 37062
rect 8186 24166 8370 36342
rect 8504 22932 8572 30498
rect 8803 21072 8871 28738
rect 8978 24166 9162 35622
rect 10674 24166 10858 35622
rect 10964 21258 11032 28738
rect 11264 23118 11332 30498
rect 11466 24166 11650 36342
rect 12042 28092 12226 37062
rect 12650 28092 12834 37062
rect 13226 24166 13410 36342
rect 13544 23304 13612 30498
rect 13843 21444 13911 28738
rect 14018 24166 14202 35622
rect 15714 24166 15898 35622
rect 16004 21630 16072 28738
rect 16304 23490 16372 30498
rect 16506 24166 16690 36342
rect 17082 28092 17266 37062
rect 17690 28092 17874 37062
rect 18266 24166 18450 36342
rect 18883 28738 18951 28922
rect 19058 24166 19242 35622
rect 20322 19856 20390 25540
rect 20598 19856 20666 30116
rect 20754 24166 20938 35622
rect 21546 24166 21730 36342
rect 8580 19516 22440 19584
rect 8580 19144 22440 19212
rect 8614 4986 10146 5054
rect 8006 -1440 8190 4800
rect 8798 -720 8982 4800
rect 9376 -1864 9444 2938
rect 10078 1178 10146 4986
rect 12210 4986 13742 5054
rect 10482 2518 12042 2586
rect 10482 1178 10550 2518
rect 12210 1178 12278 4986
rect 10078 1110 10550 1178
rect 12042 1110 12278 1178
rect 10206 230 10390 298
rect 11966 230 12150 298
rect 12912 -1864 12980 2938
rect 13374 -720 13558 4800
rect 14166 -1440 14350 4800
use SUNSAR_SARDIGEX4_CV  XA0
timestamp 1712087342
transform 1 0 -162 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARDIGEX4_CV  XA1
timestamp 1712087342
transform -1 0 4878 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARDIGEX4_CV  XA2
timestamp 1712087342
transform 1 0 4878 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARDIGEX4_CV  XA3
timestamp 1712087342
transform -1 0 9918 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARDIGEX4_CV  XA4
timestamp 1712087342
transform 1 0 9918 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARDIGEX4_CV  XA5
timestamp 1712087342
transform -1 0 14958 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARDIGEX4_CV  XA6
timestamp 1712087342
transform 1 0 14958 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARDIGEX4_CV  XA7
timestamp 1712087342
transform -1 0 19998 0 1 24166
box -180 -132 2700 10868
use SUNSAR_SARCMPX1_CV  XA20
timestamp 1712087342
transform 1 0 19998 0 1 24166
box -180 -132 2700 9988
use SUNSAR_SARBSSW_CV  XB1
timestamp 1712087342
transform -1 0 11178 0 1 0
box -180 -132 11540 4800
use SUNSAR_SARBSSW_CV  XB2
timestamp 1712087342
transform 1 0 11178 0 1 0
box -180 -132 11540 4800
use SUNSAR_cut_M3M4_1x2  xcut0
timestamp 1712008800
transform 1 0 13708 0 1 18654
box 0 0 68 184
use SUNSAR_cut_M3M4_2x1  xcut1
timestamp 1712008800
transform 1 0 13708 0 1 19144
box 0 0 184 68
use SUNSAR_cut_M3M4_1x2  xcut2
timestamp 1712008800
transform 1 0 8580 0 1 18654
box 0 0 68 184
use SUNSAR_cut_M3M4_2x1  xcut3
timestamp 1712008800
transform 1 0 8580 0 1 19516
box 0 0 184 68
use SUNSAR_cut_M2M4_2x1  xcut4
timestamp 1712008800
transform 1 0 20322 0 1 25540
box 0 0 184 68
use SUNSAR_cut_M3M4_2x1  xcut5
timestamp 1712008800
transform 1 0 20322 0 1 19516
box 0 0 184 68
use SUNSAR_cut_M3M4_1x2  xcut6
timestamp 1712008800
transform 1 0 20322 0 1 19856
box 0 0 68 184
use SUNSAR_cut_M3M4_2x1  xcut7
timestamp 1712008800
transform 1 0 20482 0 1 30116
box 0 0 184 68
use SUNSAR_cut_M2M3_2x1  xcut8
timestamp 1712008800
transform 1 0 20322 0 1 30116
box 0 0 184 68
use SUNSAR_cut_M3M4_2x1  xcut9
timestamp 1712008800
transform 1 0 20598 0 1 19144
box 0 0 184 68
use SUNSAR_cut_M3M4_1x2  xcut10
timestamp 1712008800
transform 1 0 20598 0 1 19856
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut11
timestamp 1712008800
transform 1 0 194 0 1 19830
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut12
timestamp 1712008800
transform 1 0 13156 0 1 19830
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut13
timestamp 1712008800
transform 1 0 4338 0 1 20016
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut14
timestamp 1712008800
transform 1 0 12780 0 1 20016
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut15
timestamp 1712008800
transform 1 0 5234 0 1 20202
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut16
timestamp 1712008800
transform 1 0 12404 0 1 20202
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut17
timestamp 1712008800
transform 1 0 884 0 1 20388
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut18
timestamp 1712008800
transform 1 0 9132 0 1 20388
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut19
timestamp 1712008800
transform 1 0 3763 0 1 20574
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut20
timestamp 1712008800
transform 1 0 9508 0 1 20574
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut21
timestamp 1712008800
transform 1 0 5924 0 1 20760
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut22
timestamp 1712008800
transform 1 0 9884 0 1 20760
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut23
timestamp 1712008800
transform 1 0 8803 0 1 20946
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut24
timestamp 1712008800
transform 1 0 10260 0 1 20946
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut25
timestamp 1712008800
transform 1 0 10964 0 1 21132
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut26
timestamp 1712008800
transform 1 0 10448 0 1 21132
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut27
timestamp 1712008800
transform 1 0 13843 0 1 21318
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut28
timestamp 1712008800
transform 1 0 10636 0 1 21318
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut29
timestamp 1712008800
transform 1 0 16004 0 1 21504
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut30
timestamp 1712008800
transform 1 0 10824 0 1 21504
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut31
timestamp 1712008800
transform 1 0 1027 0 1 21690
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut32
timestamp 1712008800
transform 1 0 9320 0 1 21690
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut33
timestamp 1712008800
transform 1 0 3620 0 1 21876
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut34
timestamp 1712008800
transform 1 0 9696 0 1 21876
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut35
timestamp 1712008800
transform 1 0 6067 0 1 22062
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut36
timestamp 1712008800
transform 1 0 10072 0 1 22062
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut37
timestamp 1712008800
transform 1 0 1184 0 1 22248
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut38
timestamp 1712008800
transform 1 0 12968 0 1 22248
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut39
timestamp 1712008800
transform 1 0 3464 0 1 22434
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut40
timestamp 1712008800
transform 1 0 12592 0 1 22434
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut41
timestamp 1712008800
transform 1 0 6224 0 1 22620
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut42
timestamp 1712008800
transform 1 0 12216 0 1 22620
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut43
timestamp 1712008800
transform 1 0 8504 0 1 22806
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut44
timestamp 1712008800
transform 1 0 12028 0 1 22806
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut45
timestamp 1712008800
transform 1 0 11264 0 1 22992
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut46
timestamp 1712008800
transform 1 0 11840 0 1 22992
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut47
timestamp 1712008800
transform 1 0 13544 0 1 23178
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut48
timestamp 1712008800
transform 1 0 11652 0 1 23178
box 0 0 68 184
use SUNSAR_cut_M3M4_1x2  xcut49
timestamp 1712008800
transform 1 0 16304 0 1 23364
box 0 0 68 184
use SUNSAR_cut_M2M3_1x2  xcut50
timestamp 1712008800
transform 1 0 11464 0 1 23364
box 0 0 68 184
use SUNSAR_cut_M2M4_2x2  xcut51
timestamp 1712008800
transform 1 0 594 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut52
timestamp 1712008800
transform 1 0 3938 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut53
timestamp 1712008800
transform 1 0 5634 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut54
timestamp 1712008800
transform 1 0 8978 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut55
timestamp 1712008800
transform 1 0 10674 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut56
timestamp 1712008800
transform 1 0 14018 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut57
timestamp 1712008800
transform 1 0 15714 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut58
timestamp 1712008800
transform 1 0 19058 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut59
timestamp 1712008800
transform 1 0 20754 0 1 35438
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut60
timestamp 1712008800
transform 1 0 8798 0 1 -720
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut61
timestamp 1712008800
transform 1 0 13374 0 1 -720
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut62
timestamp 1712008800
transform 1 0 1386 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut63
timestamp 1712008800
transform 1 0 3146 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut64
timestamp 1712008800
transform 1 0 6426 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut65
timestamp 1712008800
transform 1 0 8186 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut66
timestamp 1712008800
transform 1 0 11466 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut67
timestamp 1712008800
transform 1 0 13226 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut68
timestamp 1712008800
transform 1 0 16506 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut69
timestamp 1712008800
transform 1 0 18266 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut70
timestamp 1712008800
transform 1 0 21546 0 1 36158
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut71
timestamp 1712008800
transform 1 0 8006 0 1 -1440
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut72
timestamp 1712008800
transform 1 0 14166 0 1 -1440
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut73
timestamp 1712008800
transform 1 0 1962 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut74
timestamp 1712008800
transform 1 0 2570 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut75
timestamp 1712008800
transform 1 0 7002 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut76
timestamp 1712008800
transform 1 0 7610 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut77
timestamp 1712008800
transform 1 0 12042 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut78
timestamp 1712008800
transform 1 0 12650 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut79
timestamp 1712008800
transform 1 0 17082 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M2M4_2x2  xcut80
timestamp 1712008800
transform 1 0 17690 0 1 36878
box 0 0 184 184
use SUNSAR_cut_M1M3_2x1  xcut81
timestamp 1712008800
transform 1 0 9214 0 1 494
box 0 0 184 68
use SUNSAR_cut_M2M3_2x1  xcut82
timestamp 1712008800
transform 1 0 9214 0 1 -1652
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut83
timestamp 1712008800
transform 1 0 12958 0 1 494
box 0 0 184 68
use SUNSAR_cut_M2M3_2x1  xcut84
timestamp 1712008800
transform 1 0 12958 0 1 -1652
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut85
timestamp 1712008800
transform 1 0 162 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M2M3_1x2  xcut86
timestamp 1712008800
transform 1 0 -1922 0 1 33930
box 0 0 68 184
use SUNSAR_cut_M2M4_2x1  xcut87
timestamp 1712008800
transform 1 0 9318 0 1 -1864
box 0 0 184 68
use SUNSAR_cut_M2M4_2x1  xcut88
timestamp 1712008800
transform 1 0 12854 0 1 -1864
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut89
timestamp 1712008800
transform 1 0 1386 0 1 34462
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut90
timestamp 1712008800
transform 1 0 4338 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut91
timestamp 1712008800
transform 1 0 6426 0 1 34462
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut92
timestamp 1712008800
transform 1 0 9378 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut93
timestamp 1712008800
transform 1 0 11466 0 1 34462
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut94
timestamp 1712008800
transform 1 0 14418 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut95
timestamp 1712008800
transform 1 0 16506 0 1 34462
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut96
timestamp 1712008800
transform 1 0 19458 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut97
timestamp 1712008800
transform 1 0 162 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut98
timestamp 1712008800
transform 1 0 4338 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut99
timestamp 1712008800
transform 1 0 5202 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut100
timestamp 1712008800
transform 1 0 9378 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut101
timestamp 1712008800
transform 1 0 10242 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut102
timestamp 1712008800
transform 1 0 14418 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut103
timestamp 1712008800
transform 1 0 15282 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut104
timestamp 1712008800
transform 1 0 19458 0 1 31524
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut105
timestamp 1712008800
transform 1 0 3114 0 1 34428
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut106
timestamp 1712008800
transform 1 0 5202 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut107
timestamp 1712008800
transform 1 0 8154 0 1 34428
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut108
timestamp 1712008800
transform 1 0 10242 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut109
timestamp 1712008800
transform 1 0 13194 0 1 34428
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut110
timestamp 1712008800
transform 1 0 15282 0 1 33988
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut111
timestamp 1712008800
transform 1 0 162 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut112
timestamp 1712008800
transform 1 0 4338 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut113
timestamp 1712008800
transform 1 0 5202 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut114
timestamp 1712008800
transform 1 0 9378 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut115
timestamp 1712008800
transform 1 0 10242 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut116
timestamp 1712008800
transform 1 0 14418 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut117
timestamp 1712008800
transform 1 0 15282 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut118
timestamp 1712008800
transform 1 0 19458 0 1 27124
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut119
timestamp 1712008800
transform 1 0 1818 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut120
timestamp 1712008800
transform 1 0 2682 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut121
timestamp 1712008800
transform 1 0 6858 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut122
timestamp 1712008800
transform 1 0 7722 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut123
timestamp 1712008800
transform 1 0 11898 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut124
timestamp 1712008800
transform 1 0 12762 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut125
timestamp 1712008800
transform 1 0 16938 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut126
timestamp 1712008800
transform 1 0 17802 0 1 27476
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut127
timestamp 1712008800
transform 1 0 594 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut128
timestamp 1712008800
transform 1 0 3906 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut129
timestamp 1712008800
transform 1 0 5634 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut130
timestamp 1712008800
transform 1 0 8946 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut131
timestamp 1712008800
transform 1 0 10674 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut132
timestamp 1712008800
transform 1 0 13986 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut133
timestamp 1712008800
transform 1 0 15714 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut134
timestamp 1712008800
transform 1 0 19026 0 1 32668
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut135
timestamp 1712008800
transform 1 0 20322 0 1 33108
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut136
timestamp 1712008800
transform 1 0 20786 0 1 27598
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut137
timestamp 1712008800
transform 1 0 21546 0 1 28444
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut138
timestamp 1712008800
transform 1 0 21978 0 1 32932
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut139
timestamp 1712008800
transform 1 0 19458 0 1 31876
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut140
timestamp 1712008800
transform 1 0 18234 0 1 34428
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut141
timestamp 1712008800
transform 1 0 20322 0 1 33494
box 0 0 184 68
use SUNSAR_cut_M1M4_2x1  xcut142
timestamp 1712008800
transform 1 0 11934 0 1 1110
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut143
timestamp 1712008800
transform 1 0 10206 0 1 2518
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut144
timestamp 1712008800
transform 1 0 11934 0 1 1110
box 0 0 184 68
use SUNSAR_cut_M1M4_2x1  xcut145
timestamp 1712008800
transform 1 0 10206 0 1 1110
box 0 0 184 68
use SUNSAR_cut_M1M4_2x1  xcut146
timestamp 1712008800
transform 1 0 11934 0 1 2518
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut147
timestamp 1712008800
transform 1 0 162 0 1 27476
box 0 0 184 68
use SUNSAR_CDAC7_CV  XDAC1
timestamp 1712087342
transform -1 0 11028 0 1 4986
box 136 0 11028 13668
use SUNSAR_CDAC7_CV  XDAC2
timestamp 1712087342
transform 1 0 11328 0 1 4986
box 136 0 11028 13668
<< labels >>
flabel metal3 s 194 19956 262 28708 0 FreeSans 400 0 0 0 D<7>
port 6 nsew signal bidirectional
flabel metal3 s 3763 20700 3831 28738 0 FreeSans 400 0 0 0 D<6>
port 7 nsew signal bidirectional
flabel metal3 s 5924 20886 5992 28738 0 FreeSans 400 0 0 0 D<5>
port 8 nsew signal bidirectional
flabel metal3 s 8803 21072 8871 28738 0 FreeSans 400 0 0 0 D<4>
port 9 nsew signal bidirectional
flabel metal3 s 10964 21258 11032 28738 0 FreeSans 400 0 0 0 D<3>
port 10 nsew signal bidirectional
flabel metal3 s 13843 21444 13911 28738 0 FreeSans 400 0 0 0 D<2>
port 11 nsew signal bidirectional
flabel metal3 s 16004 21630 16072 28738 0 FreeSans 400 0 0 0 D<1>
port 12 nsew signal bidirectional
flabel metal1 s 23162 -720 23346 35622 0 FreeSans 400 0 0 0 AVSS
port 19 nsew signal bidirectional
flabel metal1 s 23882 -1440 24066 36342 0 FreeSans 400 0 0 0 AVDD
port 18 nsew signal bidirectional
flabel metal1 s -1710 36878 24066 37062 0 FreeSans 400 0 0 0 VREF
port 17 nsew signal bidirectional
flabel metal1 s 24210 -1652 24278 37062 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 16 nsew signal bidirectional
flabel locali s 19026 32668 19242 32736 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel metal3 s 10206 230 10390 298 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel metal3 s 11966 230 12150 298 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s 162 31524 378 31592 0 FreeSans 400 0 0 0 CK_SAMPLE
port 15 nsew signal bidirectional
flabel locali s 1818 27476 2034 27544 0 FreeSans 400 0 0 0 EN
port 14 nsew signal bidirectional
flabel locali s 10206 2518 10422 2586 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 10206 1110 10422 1178 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel metal3 s 18883 28738 18951 28922 0 FreeSans 400 0 0 0 D<0>
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -1922 -1864 24278 37062
<< end >>
