magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 1260 352
<< locali >>
rect 432 291 516 325
rect 516 291 828 325
rect 516 291 550 325
rect 1027 71 1061 281
rect 415 115 449 149
rect 415 203 449 237
rect 811 115 845 149
rect 811 203 845 237
rect 1206 66 1314 110
rect -54 66 54 110
rect 162 71 270 105
rect 990 247 1098 281
rect 162 247 270 281
rect 162 159 270 193
rect 378 291 486 325
<< m3 >>
rect 774 0 866 352
rect 378 0 470 352
rect 774 0 866 352
rect 378 0 470 352
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 88
box 0 88 630 264
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 176
box 0 176 630 352
use SUNSAR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNSAR_PCHDL MP1 
transform 1 0 630 0 1 88
box 630 88 1260 264
use SUNSAR_PCHDL MP2 
transform 1 0 630 0 1 176
box 630 176 1260 352
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 27
box 774 27 866 61
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 378 0 1 27
box 378 27 470 61
<< labels >>
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 990 247 1098 281 0 FreeSans 400 0 0 0 RST_N
port 3 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 400 0 0 0 EN
port 4 nsew signal bidirectional
flabel locali s 162 159 270 193 0 FreeSans 400 0 0 0 LCK_N
port 5 nsew signal bidirectional
flabel locali s 378 291 486 325 0 FreeSans 400 0 0 0 CHL
port 2 nsew signal bidirectional
flabel m3 s 774 0 866 352 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 378 0 470 352 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 352
<< end >>
