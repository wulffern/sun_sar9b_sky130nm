magic
tech sky130B
magscale 1 2
timestamp 1680904800
<< checkpaint >>
rect 0 0 76 200
<< m3 >>
rect 0 0 76 200
<< v3 >>
rect 6 12 70 76
rect 6 124 70 188
<< m4 >>
rect 0 0 76 200
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 76 200
<< end >>
