magic
tech sky130B
magscale 1 2
timestamp 1669849200
<< checkpaint >>
rect 0 0 200 76
<< locali >>
rect 0 0 184 68
<< viali >>
rect 12 6 68 62
rect 116 6 172 62
<< m1 >>
rect 0 0 184 68
<< v1 >>
rect 12 6 68 62
rect 116 6 172 62
<< m2 >>
rect 0 0 200 76
<< v2 >>
rect 12 6 76 70
rect 124 6 188 70
<< m3 >>
rect 0 0 200 76
<< labels >>
<< end >>
