magic
tech sky130A
timestamp 1708968222
<< locali >>
rect 378 1875 486 1909
rect 216 1831 334 1865
rect 300 1733 334 1831
rect 300 1699 550 1733
rect 516 1469 550 1699
rect 432 1435 550 1469
rect 912 1655 1044 1689
rect 216 1391 270 1425
rect 240 1357 334 1391
rect 300 985 334 1357
rect 432 995 550 1029
rect 216 951 334 985
rect 162 599 270 633
rect 300 501 334 951
rect 516 765 550 995
rect 432 731 550 765
rect 912 721 946 1655
rect 912 687 1044 721
rect 912 501 946 687
rect 300 467 432 501
rect 828 467 946 501
rect 990 423 1044 457
rect 912 389 1020 423
rect 912 325 946 389
rect 828 291 946 325
rect 162 247 270 281
<< metal1 >>
rect 828 1875 946 1909
rect 216 1655 334 1689
rect 300 1425 334 1655
rect 912 1601 946 1875
rect 912 1567 1044 1601
rect 300 1391 1162 1425
rect 912 1303 1044 1337
rect 912 1205 946 1303
rect 828 1171 946 1205
rect 216 1127 334 1161
rect 300 1029 334 1127
rect 300 995 432 1029
rect 912 897 946 1171
rect 1128 985 1162 1391
rect 1044 951 1162 985
rect 912 863 1044 897
rect 216 687 270 721
rect 240 653 334 687
rect 300 325 334 653
rect 1128 325 1162 951
rect 300 291 432 325
rect 828 291 1162 325
<< metal3 >>
rect 378 0 470 1936
rect 774 0 866 1936
use SUNSAR_TAPCELLB_CV  XA0
timestamp 1708968222
transform 1 0 0 0 1 0
box -90 -66 1350 242
use SUNSAR_IVX1_CV  XA1
timestamp 1708968222
transform 1 0 0 0 1 176
box -90 -66 1350 242
use SUNSAR_IVX1_CV  XA2
timestamp 1708968222
transform 1 0 0 0 1 352
box -90 -66 1350 242
use SUNSAR_IVTRIX1_CV  XA3
timestamp 1708968222
transform 1 0 0 0 1 528
box -90 -66 1350 330
use SUNSAR_IVTRIX1_CV  XA4
timestamp 1708968222
transform 1 0 0 0 1 792
box -90 -66 1350 330
use SUNSAR_IVX1_CV  XA5
timestamp 1708968222
transform 1 0 0 0 1 1056
box -90 -66 1350 242
use SUNSAR_IVTRIX1_CV  XA6
timestamp 1708968222
transform 1 0 0 0 1 1232
box -90 -66 1350 330
use SUNSAR_IVTRIX1_CV  XA7
timestamp 1708968222
transform 1 0 0 0 1 1496
box -90 -66 1350 330
use SUNSAR_IVX1_CV  XA8
timestamp 1708968222
transform 1 0 0 0 1 1760
box -90 -66 1350 242
use SUNSAR_cut_M1M2_2x1  xcut0
timestamp 1708902000
transform 1 0 990 0 1 951
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut1
timestamp 1708902000
transform 1 0 990 0 1 1391
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut2
timestamp 1708902000
transform 1 0 774 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut3
timestamp 1708902000
transform 1 0 162 0 1 687
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut4
timestamp 1708902000
transform 1 0 378 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut5
timestamp 1708902000
transform 1 0 162 0 1 1655
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut6
timestamp 1708902000
transform 1 0 990 0 1 1391
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut7
timestamp 1708902000
transform 1 0 162 0 1 1127
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut8
timestamp 1708902000
transform 1 0 378 0 1 995
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut9
timestamp 1708902000
transform 1 0 774 0 1 1171
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut10
timestamp 1708902000
transform 1 0 990 0 1 863
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut11
timestamp 1708902000
transform 1 0 990 0 1 1303
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut12
timestamp 1708902000
transform 1 0 774 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut13
timestamp 1708902000
transform 1 0 990 0 1 1567
box 0 0 92 34
<< labels >>
flabel locali s 162 599 270 633 0 FreeSans 200 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 200 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 378 1875 486 1909 0 FreeSans 200 0 0 0 Q
port 3 nsew signal bidirectional
flabel locali s 378 1699 486 1733 0 FreeSans 200 0 0 0 QN
port 4 nsew signal bidirectional
flabel metal3 s 774 0 866 1936 0 FreeSans 200 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel metal3 s 378 0 470 1936 0 FreeSans 200 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 1936
<< end >>
