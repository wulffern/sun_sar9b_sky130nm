magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 1260 176
<< locali >>
rect 432 115 516 149
rect 516 115 828 149
rect 516 115 550 149
rect 162 71 270 105
rect 378 115 486 149
rect 1206 66 1314 110
rect -54 66 54 110
<< poly >>
rect 162 79 1098 97
<< m3 >>
rect 774 0 866 176
rect 378 0 470 176
rect 774 0 866 176
rect 378 0 470 176
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNSAR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 27
box 774 27 866 61
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 378 0 1 27
box 378 27 470 61
<< labels >>
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 378 115 486 149 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel locali s 1206 66 1314 110 0 FreeSans 400 0 0 0 BULKP
port 3 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 BULKN
port 4 nsew signal bidirectional
flabel m3 s 774 0 866 176 0 FreeSans 400 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel m3 s 378 0 470 176 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
