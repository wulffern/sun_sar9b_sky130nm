magic
tech sky130A
magscale 1 1
timestamp 1712959200
<< checkpaint >>
rect 0 0 92 92
<< locali >>
rect 0 0 92 92
<< viali >>
rect 6 6 34 34
rect 6 58 34 86
rect 58 6 86 34
rect 58 58 86 86
<< m1 >>
rect 0 0 92 92
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 92 92
<< end >>
