magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 34 96
<< m3 >>
rect 0 0 34 92
<< v3 >>
rect 1 2 33 34
rect 1 58 33 90
<< m4 >>
rect 0 0 34 96
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 34 96
<< end >>
