magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect -826 -932 12480 18675
<< m3 >>
rect 4550 9716 11561 9750
rect 4550 9902 11561 9936
rect 10433 10088 10467 12914
rect 10571 10088 10605 15202
rect 361 10122 395 14496
rect 361 10122 395 14496
rect 2441 10215 2475 14496
rect 2881 10308 2915 14496
rect 718 10401 752 14509
rect 2145 10494 2179 14509
rect 2145 10494 2179 14509
rect 3238 10587 3272 14509
rect 3238 10587 3272 14509
rect 4665 10680 4699 14509
rect 4665 10680 4699 14509
rect 5758 10773 5792 14509
rect 5758 10773 5792 14509
rect 7185 10866 7219 14509
rect 7185 10866 7219 14509
rect 8278 10959 8312 14509
rect 8278 10959 8312 14509
rect 798 11052 832 14949
rect 2065 11145 2099 14949
rect 3318 11238 3352 14949
rect 886 11331 920 15389
rect 1978 11424 2012 15389
rect 3406 11517 3440 15389
rect 4498 11610 4532 15389
rect 5926 11703 5960 15389
rect 7018 11796 7052 15389
rect 8446 11889 8480 15389
rect 569 12227 669 17955
rect 2233 12227 2333 17955
rect 3089 12227 3189 17955
rect 4753 12227 4853 17955
rect 5609 12227 5709 17955
rect 7273 12227 7373 17955
rect 8129 12227 8229 17955
rect 9793 12227 9893 17955
rect 10649 12227 10749 17955
rect 4663 -360 4763 2400
rect 6959 -360 7059 2400
rect 965 12227 1065 18315
rect 1837 12227 1937 18315
rect 3485 12227 3585 18315
rect 4357 12227 4457 18315
rect 6005 12227 6105 18315
rect 6877 12227 6977 18315
rect 8525 12227 8625 18315
rect 9397 12227 9497 18315
rect 11045 12227 11145 18315
rect 4267 -720 4367 2400
rect 7355 -720 7455 2400
rect 1253 14190 1353 18675
rect 1549 14190 1649 18675
rect 3773 14190 3873 18675
rect 4069 14190 4169 18675
rect 6293 14190 6393 18675
rect 6589 14190 6689 18675
rect 8813 14190 8913 18675
rect 9109 14190 9209 18675
rect 4988 -932 5022 1471
rect 6700 -932 6734 1471
rect 5209 555 5429 589
rect 4569 2493 5209 2527
rect 6293 555 6479 589
rect 6479 2493 7153 2527
rect 5429 555 5513 589
rect 5513 1259 6293 1293
rect 5513 555 5547 1293
rect 5375 113 5475 151
rect 6247 113 6347 151
rect 9705 14509 9743 14609
<< m2 >>
rect 7134 9471 7168 9754
rect 4550 9471 4584 9940
rect 361 10088 6884 10122
rect 2441 10181 6696 10215
rect 2881 10274 6508 10308
rect 718 10367 4872 10401
rect 2145 10460 5060 10494
rect 3238 10553 5248 10587
rect 4665 10646 5436 10680
rect 5496 10739 5792 10773
rect 5590 10832 7219 10866
rect 5684 10925 8312 10959
rect 798 11018 4966 11052
rect 2065 11111 5154 11145
rect 3318 11204 5342 11238
rect 886 11297 6790 11331
rect 1978 11390 6602 11424
rect 3406 11483 6414 11517
rect 4498 11576 6320 11610
rect 5926 11669 6226 11703
rect 6098 11762 7052 11796
rect 6004 11855 8480 11889
rect 4908 -826 4942 281
rect 6780 -826 6814 281
rect -792 17138 353 17172
rect 965 17375 1133 17409
rect 1133 17074 2441 17108
rect 2407 17074 2441 17172
rect 1133 17074 1167 17409
rect 3485 17375 3653 17409
rect 3653 17074 4961 17108
rect 4927 17074 4961 17172
rect 3653 17074 3687 17409
rect 6005 17375 6173 17409
rect 6173 17074 7481 17108
rect 7447 17074 7481 17172
rect 6173 17074 6207 17409
rect 8525 17375 8693 17409
rect 8693 17074 10001 17108
rect 9967 17074 10001 17172
rect 8693 17074 8727 17409
rect 353 15842 10109 15876
rect 319 15842 353 15940
rect 2407 15842 2441 15940
rect 2839 15842 2873 15940
rect 4927 15842 4961 15940
rect 5359 15842 5393 15940
rect 7447 15842 7481 15940
rect 7879 15842 7913 15940
rect 9967 15842 10001 15940
rect 981 12606 1133 12640
rect 1133 12410 2441 12444
rect 2407 12410 2441 12508
rect 1133 12410 1167 12640
rect 3501 12606 3653 12640
rect 3653 12410 4961 12444
rect 4927 12410 4961 12508
rect 3653 12410 3687 12640
rect 6021 12606 6173 12640
rect 6173 12410 7481 12444
rect 7447 12410 7481 12508
rect 6173 12410 6207 12640
rect 8541 12606 8693 12640
rect 8693 12410 10001 12444
rect 9967 12410 10001 12508
rect 8693 12410 8727 12640
rect 1829 12606 1981 12640
rect 1981 12606 2015 12670
rect 1981 12670 2889 12704
rect 2855 12474 2889 12704
rect 4349 12606 4501 12640
rect 4501 12606 4535 12670
rect 4501 12670 5409 12704
rect 5375 12474 5409 12704
rect 6869 12606 7021 12640
rect 7021 12606 7055 12670
rect 7021 12670 7929 12704
rect 7895 12474 7929 12704
rect 9389 12606 9541 12640
rect 9541 12606 9575 12670
rect 369 13492 10093 13526
rect 335 13354 369 13526
rect 2407 13354 2441 13526
rect 2855 13354 2889 13526
rect 4927 13354 4961 13526
rect 5375 13354 5409 13526
rect 7447 13354 7481 13526
rect 7895 13354 7929 13526
rect 9967 13354 10001 13526
rect 353 13568 10109 13602
rect 319 13568 353 13740
rect 2407 13568 2441 13740
rect 2839 13568 2873 13740
rect 4927 13568 4961 13740
rect 5359 13568 5393 13740
rect 7447 13568 7481 13740
rect 7879 13568 7913 13740
rect 9967 13568 10001 13740
rect 461 13882 1181 13916
rect 1181 13882 1721 13916
rect 1181 13882 3809 13916
rect 1181 13882 4241 13916
rect 1181 13882 6329 13916
rect 1181 13882 6761 13916
rect 1181 13882 8849 13916
rect 1181 13882 9281 13916
rect 623 16478 707 16512
rect 707 16478 741 16512
rect 2279 16478 2363 16512
rect 2363 16478 2397 16512
rect 3143 16478 3227 16512
rect 3227 16478 3261 16512
rect 4799 16478 4883 16512
rect 4883 16478 4917 16512
rect 5663 16478 5747 16512
rect 5747 16478 5781 16512
rect 7319 16478 7403 16512
rect 7403 16478 7437 16512
rect 8183 16478 8267 16512
rect 8267 16478 8301 16512
rect 9839 16478 9923 16512
rect 9923 16698 10487 16732
rect 9923 16478 9957 16732
rect 10375 13943 10703 13977
rect 10063 13388 10375 13422
rect 10375 13388 10409 13977
rect 10047 13354 10093 13388
rect 10055 13706 10139 13740
rect 10139 14400 11075 14434
rect 10139 13706 10173 14434
rect 11045 14366 11099 14400
rect 11315 16610 11399 16644
rect 10079 16048 11399 16082
rect 11399 16048 11433 16644
rect 10055 16082 10109 16116
rect 9443 17358 10205 17392
rect 10205 16891 10487 16925
rect 10205 16891 10239 17392
rect 5429 1259 5513 1293
rect 5513 555 6293 589
rect 5513 555 5547 1293
rect 353 13882 1289 13916
<< m4 >>
rect 10433 9902 10467 10088
rect 10571 9716 10605 10088
rect 5209 555 5243 2527
rect 6479 555 6513 2527
<< m1 >>
rect 6850 9437 6884 10088
rect 6662 9437 6696 10181
rect 6474 9437 6508 10274
rect 4838 9437 4872 10367
rect 5026 9437 5060 10460
rect 5214 9437 5248 10553
rect 5402 9437 5436 10646
rect 5496 9437 5530 10739
rect 5590 9437 5624 10832
rect 5684 9437 5718 10925
rect 4932 9437 4966 11018
rect 5120 9437 5154 11111
rect 5308 9437 5342 11204
rect 6756 9437 6790 11297
rect 6568 9437 6602 11390
rect 6380 9437 6414 11483
rect 6286 9437 6320 11576
rect 6192 9437 6226 11669
rect 6098 9437 6132 11762
rect 6004 9437 6038 11855
rect 11914 -360 12014 17955
rect -360 -360 12014 -260
rect -360 17855 12014 17955
rect -360 -360 -260 17955
rect 11914 -360 12014 17955
rect 12274 -720 12374 18315
rect -720 -720 12374 -620
rect -720 18215 12374 18315
rect -720 -720 -620 18315
rect 12274 -720 12374 18315
rect -720 18575 12374 18675
rect -720 18575 12374 18675
rect 12446 -826 12480 18675
rect -720 -826 12480 -792
rect 12446 -826 12480 18675
rect -826 -932 12480 -898
rect -826 -932 -792 18675
rect 1829 17358 1997 17392
rect 1997 17074 2873 17108
rect 2839 17074 2873 17172
rect 1997 17074 2031 17392
rect 4349 17358 4517 17392
rect 4517 17074 5393 17108
rect 5359 17074 5393 17172
rect 4517 17074 4551 17392
rect 6869 17358 7037 17392
rect 7037 17074 7913 17108
rect 7879 17074 7913 17172
rect 7037 17074 7071 17392
rect -360 2493 38 2527
rect -360 4229 38 4263
rect -360 5965 38 5999
rect -360 7701 38 7735
rect 11684 2493 12014 2527
rect 11684 4229 12014 4263
rect 11684 5965 12014 5999
rect 11684 7701 12014 7735
<< locali >>
rect 9785 16478 9893 16512
rect 353 15906 461 15940
rect 1181 13882 1289 13916
rect 5375 1259 5483 1293
rect 5375 555 5483 589
use SUNSAR_SARBSSW_CV XB1 
transform -1 0 5861 0 1 0
box 5861 0 11585 2400
use SUNSAR_SARBSSW_CV XB2 
transform 1 0 5861 0 1 0
box 5861 0 11585 2400
use SUNSAR_CDAC7_CV XDAC1 
transform -1 0 5786 0 1 2493
box 5786 2493 11504 9471
use SUNSAR_CDAC7_CV XDAC2 
transform 1 0 5936 0 1 2493
box 5936 2493 11654 9471
use SUNSAR_SARDIGEX4_CV XA0 
transform 1 0 191 0 1 12227
box 191 12227 1451 17595
use SUNSAR_SARDIGEX4_CV XA1 
transform -1 0 2711 0 1 12227
box 2711 12227 3971 17595
use SUNSAR_SARDIGEX4_CV XA2 
transform 1 0 2711 0 1 12227
box 2711 12227 3971 17595
use SUNSAR_SARDIGEX4_CV XA3 
transform -1 0 5231 0 1 12227
box 5231 12227 6491 17595
use SUNSAR_SARDIGEX4_CV XA4 
transform 1 0 5231 0 1 12227
box 5231 12227 6491 17595
use SUNSAR_SARDIGEX4_CV XA5 
transform -1 0 7751 0 1 12227
box 7751 12227 9011 17595
use SUNSAR_SARDIGEX4_CV XA6 
transform 1 0 7751 0 1 12227
box 7751 12227 9011 17595
use SUNSAR_SARDIGEX4_CV XA7 
transform -1 0 10271 0 1 12227
box 10271 12227 11531 17595
use SUNSAR_SARCMPX1_CV XA20 
transform 1 0 10271 0 1 12227
box 10271 12227 11531 17155
use SUNSAR_cut_M3M4_1x2 xcut0 
transform 1 0 7134 0 1 9471
box 7134 9471 7172 9571
use SUNSAR_cut_M3M4_2x1 xcut1 
transform 1 0 7134 0 1 9716
box 7134 9716 7234 9754
use SUNSAR_cut_M3M4_1x2 xcut2 
transform 1 0 4550 0 1 9471
box 4550 9471 4588 9571
use SUNSAR_cut_M3M4_2x1 xcut3 
transform 1 0 4550 0 1 9902
box 4550 9902 4650 9940
use SUNSAR_cut_M2M4_2x1 xcut4 
transform 1 0 10433 0 1 12914
box 10433 12914 10533 12952
use SUNSAR_cut_M4M5_2x1 xcut5 
transform 1 0 10433 0 1 9902
box 10433 9902 10533 9940
use SUNSAR_cut_M4M5_1x2 xcut6 
transform 1 0 10433 0 1 10088
box 10433 10088 10471 10188
use SUNSAR_cut_M3M4_2x1 xcut7 
transform 1 0 10513 0 1 15202
box 10513 15202 10613 15240
use SUNSAR_cut_M2M3_2x1 xcut8 
transform 1 0 10433 0 1 15202
box 10433 15202 10525 15236
use SUNSAR_cut_M4M5_2x1 xcut9 
transform 1 0 10571 0 1 9716
box 10571 9716 10671 9754
use SUNSAR_cut_M4M5_1x2 xcut10 
transform 1 0 10571 0 1 10088
box 10571 10088 10609 10188
use SUNSAR_cut_M3M4_1x2 xcut11 
transform 1 0 359 0 1 10055
box 359 10055 397 10155
use SUNSAR_cut_M2M3_1x2 xcut12 
transform 1 0 6850 0 1 10059
box 6850 10059 6884 10151
use SUNSAR_cut_M3M4_1x2 xcut13 
transform 1 0 2439 0 1 10148
box 2439 10148 2477 10248
use SUNSAR_cut_M2M3_1x2 xcut14 
transform 1 0 6662 0 1 10152
box 6662 10152 6696 10244
use SUNSAR_cut_M3M4_1x2 xcut15 
transform 1 0 2879 0 1 10241
box 2879 10241 2917 10341
use SUNSAR_cut_M2M3_1x2 xcut16 
transform 1 0 6474 0 1 10245
box 6474 10245 6508 10337
use SUNSAR_cut_M3M4_1x2 xcut17 
transform 1 0 716 0 1 10334
box 716 10334 754 10434
use SUNSAR_cut_M2M3_1x2 xcut18 
transform 1 0 4838 0 1 10338
box 4838 10338 4872 10430
use SUNSAR_cut_M3M4_1x2 xcut19 
transform 1 0 2143 0 1 10427
box 2143 10427 2181 10527
use SUNSAR_cut_M2M3_1x2 xcut20 
transform 1 0 5026 0 1 10431
box 5026 10431 5060 10523
use SUNSAR_cut_M3M4_1x2 xcut21 
transform 1 0 3236 0 1 10520
box 3236 10520 3274 10620
use SUNSAR_cut_M2M3_1x2 xcut22 
transform 1 0 5214 0 1 10524
box 5214 10524 5248 10616
use SUNSAR_cut_M3M4_1x2 xcut23 
transform 1 0 4663 0 1 10613
box 4663 10613 4701 10713
use SUNSAR_cut_M2M3_1x2 xcut24 
transform 1 0 5402 0 1 10617
box 5402 10617 5436 10709
use SUNSAR_cut_M3M4_1x2 xcut25 
transform 1 0 5756 0 1 10706
box 5756 10706 5794 10806
use SUNSAR_cut_M2M3_1x2 xcut26 
transform 1 0 5496 0 1 10710
box 5496 10710 5530 10802
use SUNSAR_cut_M3M4_1x2 xcut27 
transform 1 0 7183 0 1 10799
box 7183 10799 7221 10899
use SUNSAR_cut_M2M3_1x2 xcut28 
transform 1 0 5590 0 1 10803
box 5590 10803 5624 10895
use SUNSAR_cut_M3M4_1x2 xcut29 
transform 1 0 8276 0 1 10892
box 8276 10892 8314 10992
use SUNSAR_cut_M2M3_1x2 xcut30 
transform 1 0 5684 0 1 10896
box 5684 10896 5718 10988
use SUNSAR_cut_M3M4_1x2 xcut31 
transform 1 0 796 0 1 10985
box 796 10985 834 11085
use SUNSAR_cut_M2M3_1x2 xcut32 
transform 1 0 4932 0 1 10989
box 4932 10989 4966 11081
use SUNSAR_cut_M3M4_1x2 xcut33 
transform 1 0 2063 0 1 11078
box 2063 11078 2101 11178
use SUNSAR_cut_M2M3_1x2 xcut34 
transform 1 0 5120 0 1 11082
box 5120 11082 5154 11174
use SUNSAR_cut_M3M4_1x2 xcut35 
transform 1 0 3316 0 1 11171
box 3316 11171 3354 11271
use SUNSAR_cut_M2M3_1x2 xcut36 
transform 1 0 5308 0 1 11175
box 5308 11175 5342 11267
use SUNSAR_cut_M3M4_1x2 xcut37 
transform 1 0 884 0 1 11264
box 884 11264 922 11364
use SUNSAR_cut_M2M3_1x2 xcut38 
transform 1 0 6756 0 1 11268
box 6756 11268 6790 11360
use SUNSAR_cut_M3M4_1x2 xcut39 
transform 1 0 1976 0 1 11357
box 1976 11357 2014 11457
use SUNSAR_cut_M2M3_1x2 xcut40 
transform 1 0 6568 0 1 11361
box 6568 11361 6602 11453
use SUNSAR_cut_M3M4_1x2 xcut41 
transform 1 0 3404 0 1 11450
box 3404 11450 3442 11550
use SUNSAR_cut_M2M3_1x2 xcut42 
transform 1 0 6380 0 1 11454
box 6380 11454 6414 11546
use SUNSAR_cut_M3M4_1x2 xcut43 
transform 1 0 4496 0 1 11543
box 4496 11543 4534 11643
use SUNSAR_cut_M2M3_1x2 xcut44 
transform 1 0 6286 0 1 11547
box 6286 11547 6320 11639
use SUNSAR_cut_M3M4_1x2 xcut45 
transform 1 0 5924 0 1 11636
box 5924 11636 5962 11736
use SUNSAR_cut_M2M3_1x2 xcut46 
transform 1 0 6192 0 1 11640
box 6192 11640 6226 11732
use SUNSAR_cut_M3M4_1x2 xcut47 
transform 1 0 7016 0 1 11729
box 7016 11729 7054 11829
use SUNSAR_cut_M2M3_1x2 xcut48 
transform 1 0 6098 0 1 11733
box 6098 11733 6132 11825
use SUNSAR_cut_M3M4_1x2 xcut49 
transform 1 0 8444 0 1 11822
box 8444 11822 8482 11922
use SUNSAR_cut_M2M3_1x2 xcut50 
transform 1 0 6004 0 1 11826
box 6004 11826 6038 11918
use SUNSAR_cut_M2M4_2x2 xcut51 
transform 1 0 569 0 1 17855
box 569 17855 669 17955
use SUNSAR_cut_M2M4_2x2 xcut52 
transform 1 0 2233 0 1 17855
box 2233 17855 2333 17955
use SUNSAR_cut_M2M4_2x2 xcut53 
transform 1 0 3089 0 1 17855
box 3089 17855 3189 17955
use SUNSAR_cut_M2M4_2x2 xcut54 
transform 1 0 4753 0 1 17855
box 4753 17855 4853 17955
use SUNSAR_cut_M2M4_2x2 xcut55 
transform 1 0 5609 0 1 17855
box 5609 17855 5709 17955
use SUNSAR_cut_M2M4_2x2 xcut56 
transform 1 0 7273 0 1 17855
box 7273 17855 7373 17955
use SUNSAR_cut_M2M4_2x2 xcut57 
transform 1 0 8129 0 1 17855
box 8129 17855 8229 17955
use SUNSAR_cut_M2M4_2x2 xcut58 
transform 1 0 9793 0 1 17855
box 9793 17855 9893 17955
use SUNSAR_cut_M2M4_2x2 xcut59 
transform 1 0 10649 0 1 17855
box 10649 17855 10749 17955
use SUNSAR_cut_M2M4_2x2 xcut60 
transform 1 0 4663 0 1 -360
box 4663 -360 4763 -260
use SUNSAR_cut_M2M4_2x2 xcut61 
transform 1 0 6959 0 1 -360
box 6959 -360 7059 -260
use SUNSAR_cut_M2M4_2x2 xcut62 
transform 1 0 965 0 1 18215
box 965 18215 1065 18315
use SUNSAR_cut_M2M4_2x2 xcut63 
transform 1 0 1837 0 1 18215
box 1837 18215 1937 18315
use SUNSAR_cut_M2M4_2x2 xcut64 
transform 1 0 3485 0 1 18215
box 3485 18215 3585 18315
use SUNSAR_cut_M2M4_2x2 xcut65 
transform 1 0 4357 0 1 18215
box 4357 18215 4457 18315
use SUNSAR_cut_M2M4_2x2 xcut66 
transform 1 0 6005 0 1 18215
box 6005 18215 6105 18315
use SUNSAR_cut_M2M4_2x2 xcut67 
transform 1 0 6877 0 1 18215
box 6877 18215 6977 18315
use SUNSAR_cut_M2M4_2x2 xcut68 
transform 1 0 8525 0 1 18215
box 8525 18215 8625 18315
use SUNSAR_cut_M2M4_2x2 xcut69 
transform 1 0 9397 0 1 18215
box 9397 18215 9497 18315
use SUNSAR_cut_M2M4_2x2 xcut70 
transform 1 0 11045 0 1 18215
box 11045 18215 11145 18315
use SUNSAR_cut_M2M4_2x2 xcut71 
transform 1 0 4267 0 1 -720
box 4267 -720 4367 -620
use SUNSAR_cut_M2M4_2x2 xcut72 
transform 1 0 7355 0 1 -720
box 7355 -720 7455 -620
use SUNSAR_cut_M2M4_2x2 xcut73 
transform 1 0 1253 0 1 18575
box 1253 18575 1353 18675
use SUNSAR_cut_M2M4_2x2 xcut74 
transform 1 0 1549 0 1 18575
box 1549 18575 1649 18675
use SUNSAR_cut_M2M4_2x2 xcut75 
transform 1 0 3773 0 1 18575
box 3773 18575 3873 18675
use SUNSAR_cut_M2M4_2x2 xcut76 
transform 1 0 4069 0 1 18575
box 4069 18575 4169 18675
use SUNSAR_cut_M2M4_2x2 xcut77 
transform 1 0 6293 0 1 18575
box 6293 18575 6393 18675
use SUNSAR_cut_M2M4_2x2 xcut78 
transform 1 0 6589 0 1 18575
box 6589 18575 6689 18675
use SUNSAR_cut_M2M4_2x2 xcut79 
transform 1 0 8813 0 1 18575
box 8813 18575 8913 18675
use SUNSAR_cut_M2M4_2x2 xcut80 
transform 1 0 9109 0 1 18575
box 9109 18575 9209 18675
use SUNSAR_cut_M1M3_2x1 xcut81 
transform 1 0 4879 0 1 247
box 4879 247 4971 281
use SUNSAR_cut_M2M3_2x1 xcut82 
transform 1 0 4879 0 1 -826
box 4879 -826 4971 -792
use SUNSAR_cut_M1M3_2x1 xcut83 
transform 1 0 6751 0 1 247
box 6751 247 6843 281
use SUNSAR_cut_M2M3_2x1 xcut84 
transform 1 0 6751 0 1 -826
box 6751 -826 6843 -792
use SUNSAR_cut_M1M3_2x1 xcut85 
transform 1 0 353 0 1 17138
box 353 17138 445 17172
use SUNSAR_cut_M2M3_1x2 xcut86 
transform 1 0 -826 0 1 17109
box -826 17109 -792 17201
use SUNSAR_cut_M2M4_2x1 xcut87 
transform 1 0 4955 0 1 -932
box 4955 -932 5055 -894
use SUNSAR_cut_M2M4_2x1 xcut88 
transform 1 0 6667 0 1 -932
box 6667 -932 6767 -894
use SUNSAR_cut_M1M3_2x1 xcut89 
transform 1 0 965 0 1 17375
box 965 17375 1057 17409
use SUNSAR_cut_M1M3_2x1 xcut90 
transform 1 0 2441 0 1 17138
box 2441 17138 2533 17172
use SUNSAR_cut_M1M3_2x1 xcut91 
transform 1 0 3485 0 1 17375
box 3485 17375 3577 17409
use SUNSAR_cut_M1M3_2x1 xcut92 
transform 1 0 4961 0 1 17138
box 4961 17138 5053 17172
use SUNSAR_cut_M1M3_2x1 xcut93 
transform 1 0 6005 0 1 17375
box 6005 17375 6097 17409
use SUNSAR_cut_M1M3_2x1 xcut94 
transform 1 0 7481 0 1 17138
box 7481 17138 7573 17172
use SUNSAR_cut_M1M3_2x1 xcut95 
transform 1 0 8525 0 1 17375
box 8525 17375 8617 17409
use SUNSAR_cut_M1M3_2x1 xcut96 
transform 1 0 10001 0 1 17138
box 10001 17138 10093 17172
use SUNSAR_cut_M1M3_2x1 xcut97 
transform 1 0 353 0 1 15906
box 353 15906 445 15940
use SUNSAR_cut_M1M3_2x1 xcut98 
transform 1 0 2441 0 1 15906
box 2441 15906 2533 15940
use SUNSAR_cut_M1M3_2x1 xcut99 
transform 1 0 2873 0 1 15906
box 2873 15906 2965 15940
use SUNSAR_cut_M1M3_2x1 xcut100 
transform 1 0 4961 0 1 15906
box 4961 15906 5053 15940
use SUNSAR_cut_M1M3_2x1 xcut101 
transform 1 0 5393 0 1 15906
box 5393 15906 5485 15940
use SUNSAR_cut_M1M3_2x1 xcut102 
transform 1 0 7481 0 1 15906
box 7481 15906 7573 15940
use SUNSAR_cut_M1M3_2x1 xcut103 
transform 1 0 7913 0 1 15906
box 7913 15906 8005 15940
use SUNSAR_cut_M1M3_2x1 xcut104 
transform 1 0 10001 0 1 15906
box 10001 15906 10093 15940
use SUNSAR_cut_M1M2_2x1 xcut105 
transform 1 0 1829 0 1 17358
box 1829 17358 1921 17392
use SUNSAR_cut_M1M2_2x1 xcut106 
transform 1 0 2873 0 1 17138
box 2873 17138 2965 17172
use SUNSAR_cut_M1M2_2x1 xcut107 
transform 1 0 4349 0 1 17358
box 4349 17358 4441 17392
use SUNSAR_cut_M1M2_2x1 xcut108 
transform 1 0 5393 0 1 17138
box 5393 17138 5485 17172
use SUNSAR_cut_M1M2_2x1 xcut109 
transform 1 0 6869 0 1 17358
box 6869 17358 6961 17392
use SUNSAR_cut_M1M2_2x1 xcut110 
transform 1 0 7913 0 1 17138
box 7913 17138 8005 17172
use SUNSAR_cut_M1M3_2x1 xcut111 
transform 1 0 353 0 1 13706
box 353 13706 445 13740
use SUNSAR_cut_M1M3_2x1 xcut112 
transform 1 0 2441 0 1 13706
box 2441 13706 2533 13740
use SUNSAR_cut_M1M3_2x1 xcut113 
transform 1 0 2873 0 1 13706
box 2873 13706 2965 13740
use SUNSAR_cut_M1M3_2x1 xcut114 
transform 1 0 4961 0 1 13706
box 4961 13706 5053 13740
use SUNSAR_cut_M1M3_2x1 xcut115 
transform 1 0 5393 0 1 13706
box 5393 13706 5485 13740
use SUNSAR_cut_M1M3_2x1 xcut116 
transform 1 0 7481 0 1 13706
box 7481 13706 7573 13740
use SUNSAR_cut_M1M3_2x1 xcut117 
transform 1 0 7913 0 1 13706
box 7913 13706 8005 13740
use SUNSAR_cut_M1M3_2x1 xcut118 
transform 1 0 10001 0 1 13706
box 10001 13706 10093 13740
use SUNSAR_cut_M1M3_2x1 xcut119 
transform 1 0 1181 0 1 13882
box 1181 13882 1273 13916
use SUNSAR_cut_M1M3_2x1 xcut120 
transform 1 0 1613 0 1 13882
box 1613 13882 1705 13916
use SUNSAR_cut_M1M3_2x1 xcut121 
transform 1 0 3701 0 1 13882
box 3701 13882 3793 13916
use SUNSAR_cut_M1M3_2x1 xcut122 
transform 1 0 4133 0 1 13882
box 4133 13882 4225 13916
use SUNSAR_cut_M1M3_2x1 xcut123 
transform 1 0 6221 0 1 13882
box 6221 13882 6313 13916
use SUNSAR_cut_M1M3_2x1 xcut124 
transform 1 0 6653 0 1 13882
box 6653 13882 6745 13916
use SUNSAR_cut_M1M3_2x1 xcut125 
transform 1 0 8741 0 1 13882
box 8741 13882 8833 13916
use SUNSAR_cut_M1M3_2x1 xcut126 
transform 1 0 9173 0 1 13882
box 9173 13882 9265 13916
use SUNSAR_cut_M1M3_2x1 xcut127 
transform 1 0 569 0 1 16478
box 569 16478 661 16512
use SUNSAR_cut_M1M3_2x1 xcut128 
transform 1 0 2225 0 1 16478
box 2225 16478 2317 16512
use SUNSAR_cut_M1M3_2x1 xcut129 
transform 1 0 3089 0 1 16478
box 3089 16478 3181 16512
use SUNSAR_cut_M1M3_2x1 xcut130 
transform 1 0 4745 0 1 16478
box 4745 16478 4837 16512
use SUNSAR_cut_M1M3_2x1 xcut131 
transform 1 0 5609 0 1 16478
box 5609 16478 5701 16512
use SUNSAR_cut_M1M3_2x1 xcut132 
transform 1 0 7265 0 1 16478
box 7265 16478 7357 16512
use SUNSAR_cut_M1M3_2x1 xcut133 
transform 1 0 8129 0 1 16478
box 8129 16478 8221 16512
use SUNSAR_cut_M1M3_2x1 xcut134 
transform 1 0 9785 0 1 16478
box 9785 16478 9877 16512
use SUNSAR_cut_M1M3_2x1 xcut135 
transform 1 0 10433 0 1 16698
box 10433 16698 10525 16732
use SUNSAR_cut_M1M3_2x1 xcut136 
transform 1 0 10665 0 1 13943
box 10665 13943 10757 13977
use SUNSAR_cut_M1M3_2x1 xcut137 
transform 1 0 11045 0 1 14366
box 11045 14366 11137 14400
use SUNSAR_cut_M1M3_2x1 xcut138 
transform 1 0 11261 0 1 16610
box 11261 16610 11353 16644
use SUNSAR_cut_M1M3_2x1 xcut139 
transform 1 0 10001 0 1 16082
box 10001 16082 10093 16116
use SUNSAR_cut_M1M3_2x1 xcut140 
transform 1 0 9389 0 1 17358
box 9389 17358 9481 17392
use SUNSAR_cut_M1M3_2x1 xcut141 
transform 1 0 10433 0 1 16891
box 10433 16891 10525 16925
use SUNSAR_cut_M4M5_1x2 xcut142 
transform 1 0 5209 0 1 555
box 5209 555 5247 655
use SUNSAR_cut_M4M5_1x2 xcut143 
transform 1 0 5209 0 1 2427
box 5209 2427 5247 2527
use SUNSAR_cut_M1M4_2x1 xcut144 
transform 1 0 6239 0 1 555
box 6239 555 6339 593
use SUNSAR_cut_M4M5_1x2 xcut145 
transform 1 0 6479 0 1 555
box 6479 555 6517 655
use SUNSAR_cut_M4M5_1x2 xcut146 
transform 1 0 6479 0 1 2427
box 6479 2427 6517 2527
use SUNSAR_cut_M1M3_2x1 xcut147 
transform 1 0 5375 0 1 1259
box 5375 1259 5467 1293
use SUNSAR_cut_M1M3_2x1 xcut148 
transform 1 0 6239 0 1 555
box 6239 555 6331 589
use SUNSAR_cut_M1M4_2x1 xcut149 
transform 1 0 5375 0 1 555
box 5375 555 5475 593
use SUNSAR_cut_M1M4_2x1 xcut150 
transform 1 0 6239 0 1 1259
box 6239 1259 6339 1297
use SUNSAR_cut_M1M3_2x1 xcut151 
transform 1 0 353 0 1 13882
box 353 13882 445 13916
<< labels >>
flabel m3 s 361 10122 395 14496 0 FreeSans 400 0 0 0 D<7>
port 6 nsew signal bidirectional
flabel m3 s 2145 10494 2179 14509 0 FreeSans 400 0 0 0 D<6>
port 7 nsew signal bidirectional
flabel m3 s 3238 10587 3272 14509 0 FreeSans 400 0 0 0 D<5>
port 8 nsew signal bidirectional
flabel m3 s 4665 10680 4699 14509 0 FreeSans 400 0 0 0 D<4>
port 9 nsew signal bidirectional
flabel m3 s 5758 10773 5792 14509 0 FreeSans 400 0 0 0 D<3>
port 10 nsew signal bidirectional
flabel m3 s 7185 10866 7219 14509 0 FreeSans 400 0 0 0 D<2>
port 11 nsew signal bidirectional
flabel m3 s 8278 10959 8312 14509 0 FreeSans 400 0 0 0 D<1>
port 12 nsew signal bidirectional
flabel m1 s 11914 -360 12014 17955 0 FreeSans 400 0 0 0 AVSS
port 19 nsew signal bidirectional
flabel m1 s 12274 -720 12374 18315 0 FreeSans 400 0 0 0 AVDD
port 18 nsew signal bidirectional
flabel m1 s -720 18575 12374 18675 0 FreeSans 400 0 0 0 VREF
port 17 nsew signal bidirectional
flabel m1 s 12446 -826 12480 18675 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 16 nsew signal bidirectional
flabel locali s 9785 16478 9893 16512 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel m3 s 5375 113 5475 151 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel m3 s 6247 113 6347 151 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s 353 15906 461 15940 0 FreeSans 400 0 0 0 CK_SAMPLE
port 15 nsew signal bidirectional
flabel locali s 1181 13882 1289 13916 0 FreeSans 400 0 0 0 EN
port 14 nsew signal bidirectional
flabel locali s 5375 1259 5483 1293 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 5375 555 5483 589 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel m3 s 9705 14509 9743 14609 0 FreeSans 400 0 0 0 D<0>
port 13 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -826 -932 12480 18675
<< end >>
