magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect -1349 -932 12903 25703
<< m3 >>
rect 4290 16372 11984 16406
rect 4290 16558 11984 16592
rect 11807 16728 11841 19942
rect 11945 16728 11979 22230
rect -345 16778 -311 21526
rect -345 16778 -311 21526
rect 4247 16871 4281 21526
rect 2175 16964 2209 21526
rect 1727 17057 1761 21526
rect 0 17150 34 21541
rect 3959 17243 3993 21541
rect 3959 17243 3993 21541
rect 5040 17336 5074 21541
rect 5040 17336 5074 21541
rect 6479 17429 6513 21541
rect 6479 17429 6513 21541
rect 7560 17522 7594 21541
rect 7560 17522 7594 21541
rect 8999 17615 9033 21541
rect 8999 17615 9033 21541
rect 2520 17708 2554 21541
rect 2520 17708 2554 21541
rect 1439 17801 1473 21541
rect 1439 17801 1473 21541
rect 2591 17894 2625 21981
rect 3888 17987 3922 21981
rect 1368 18080 1402 21981
rect 71 18173 105 21981
rect 150 18266 184 22421
rect 1290 18359 1324 22421
rect 2670 18452 2704 22421
rect 3810 18545 3844 22421
rect 5190 18638 5224 22421
rect 6330 18731 6364 22421
rect 7710 18824 7744 22421
rect 8850 18917 8884 22421
rect -145 19255 -53 24983
rect 1527 19255 1619 24983
rect 2375 19255 2467 24983
rect 4047 19255 4139 24983
rect 4895 19255 4987 24983
rect 6567 19255 6659 24983
rect 7415 19255 7507 24983
rect 9087 19255 9179 24983
rect 9935 19255 10027 24983
rect 11607 19255 11699 24983
rect 4587 -360 4679 2400
rect 6875 -360 6967 2400
rect 251 19255 343 25343
rect 1131 19255 1223 25343
rect 2771 19255 2863 25343
rect 3651 19255 3743 25343
rect 5291 19255 5383 25343
rect 6171 19255 6263 25343
rect 7811 19255 7903 25343
rect 8691 19255 8783 25343
rect 10331 19255 10423 25343
rect 11211 19255 11303 25343
rect 4191 -720 4283 2400
rect 7271 -720 7363 2400
rect 539 21218 631 25703
rect 843 21218 935 25703
rect 3059 21218 3151 25703
rect 3363 21218 3455 25703
rect 5579 21218 5671 25703
rect 5883 21218 5975 25703
rect 8099 21218 8191 25703
rect 8403 21218 8495 25703
rect 10619 21218 10711 25703
rect 4876 -932 4910 1469
rect 6644 -932 6678 1469
rect 5227 555 5345 589
rect 4307 2493 5227 2527
rect 6209 555 6293 589
rect 6293 2493 7247 2527
rect 5345 555 5429 589
rect 5429 1259 6209 1293
rect 5429 555 5463 1293
rect 5291 115 5383 149
rect 6171 115 6263 149
rect 10080 21541 10114 21633
<< m2 >>
rect 7230 16127 7264 16406
rect 4290 16127 4324 16592
rect -345 16744 6988 16778
rect 4247 16837 6424 16871
rect 2175 16930 6612 16964
rect 1727 17023 6800 17057
rect 0 17116 4600 17150
rect 3959 17209 5164 17243
rect 5040 17302 5352 17336
rect 5412 17395 6513 17429
rect 5506 17488 7594 17522
rect 5600 17581 9033 17615
rect 2520 17674 4976 17708
rect 1439 17767 4788 17801
rect 2591 17860 5070 17894
rect 3888 17953 5258 17987
rect 1368 18046 4882 18080
rect 71 18139 4694 18173
rect 150 18232 6894 18266
rect 1290 18325 6706 18359
rect 2670 18418 6518 18452
rect 3810 18511 6330 18545
rect 5190 18604 6236 18638
rect 6108 18697 6364 18731
rect 6014 18790 7744 18824
rect 5920 18883 8884 18917
rect 251 24403 419 24437
rect 419 24102 1727 24136
rect 1693 24102 1727 24200
rect 419 24102 453 24437
rect 2771 24403 2939 24437
rect 2939 24102 4247 24136
rect 4213 24102 4247 24200
rect 2939 24102 2973 24437
rect 5291 24403 5459 24437
rect 5459 24102 6767 24136
rect 6733 24102 6767 24200
rect 5459 24102 5493 24437
rect 7811 24403 7979 24437
rect 7979 24102 9287 24136
rect 9253 24102 9287 24200
rect 7979 24102 8013 24437
rect -361 22870 9827 22904
rect -395 22870 -361 22968
rect 1693 22870 1727 22968
rect 2125 22870 2159 22968
rect 4213 22870 4247 22968
rect 4645 22870 4679 22968
rect 6733 22870 6767 22968
rect 7165 22870 7199 22968
rect 9253 22870 9287 22968
rect 9685 22870 9719 22968
rect 267 19634 419 19668
rect 419 19438 1727 19472
rect 1693 19438 1727 19536
rect 419 19438 453 19668
rect 2787 19634 2939 19668
rect 2939 19438 4247 19472
rect 4213 19438 4247 19536
rect 2939 19438 2973 19668
rect 5307 19634 5459 19668
rect 5459 19438 6767 19472
rect 6733 19438 6767 19536
rect 5459 19438 5493 19668
rect 7827 19634 7979 19668
rect 7979 19438 9287 19472
rect 9253 19438 9287 19536
rect 7979 19438 8013 19668
rect 10347 19634 10499 19668
rect 10499 19634 10533 19668
rect 1115 19634 1267 19668
rect 1267 19634 1301 19698
rect 1267 19698 2175 19732
rect 2141 19502 2175 19732
rect 3635 19634 3787 19668
rect 3787 19634 3821 19698
rect 3787 19698 4695 19732
rect 4661 19502 4695 19732
rect 6155 19634 6307 19668
rect 6307 19634 6341 19698
rect 6307 19698 7215 19732
rect 7181 19502 7215 19732
rect 8675 19634 8827 19668
rect 8827 19634 8861 19698
rect 8827 19698 9735 19732
rect 9701 19502 9735 19732
rect -345 20520 9827 20554
rect -379 20382 -345 20554
rect 1693 20382 1727 20554
rect 2141 20382 2175 20554
rect 4213 20382 4247 20554
rect 4661 20382 4695 20554
rect 6733 20382 6767 20554
rect 7181 20382 7215 20554
rect 9253 20382 9287 20554
rect 9701 20382 9735 20554
rect -361 20596 9827 20630
rect -395 20596 -361 20768
rect 1693 20596 1727 20768
rect 2125 20596 2159 20768
rect 4213 20596 4247 20768
rect 4645 20596 4679 20768
rect 6733 20596 6767 20768
rect 7165 20596 7199 20768
rect 9253 20596 9287 20768
rect 9685 20596 9719 20768
rect -253 20910 467 20944
rect 467 20910 1007 20944
rect 467 20910 3095 20944
rect 467 20910 3527 20944
rect 467 20910 5615 20944
rect 467 20910 6047 20944
rect 467 20910 8135 20944
rect 467 20910 8567 20944
rect 467 20910 10655 20944
rect 11461 20971 11645 21005
rect 9797 20416 11461 20450
rect 11461 20416 11495 21005
rect 9781 20382 9827 20416
rect 11131 21411 11249 21445
rect 9797 20768 11131 20802
rect 11131 20768 11165 21445
rect 9773 20734 9827 20768
rect 11033 23638 11117 23672
rect 9773 23110 11117 23144
rect 11117 23110 11151 23672
rect 10915 23902 11033 23936
rect 10385 24403 10915 24437
rect 10915 23902 10949 24437
rect 5345 1259 5429 1293
rect 5429 555 6209 589
rect 5429 555 5463 1293
rect -361 20910 575 20944
<< m4 >>
rect 11807 16558 11841 16728
rect 11945 16372 11979 16728
rect 5227 555 5261 2527
rect 6293 555 6327 2527
<< m1 >>
rect 6954 16093 6988 16744
rect 6390 16093 6424 16837
rect 6578 16093 6612 16930
rect 6766 16093 6800 17023
rect 4566 16093 4600 17116
rect 5130 16093 5164 17209
rect 5318 16093 5352 17302
rect 5412 16093 5446 17395
rect 5506 16093 5540 17488
rect 5600 16093 5634 17581
rect 4942 16093 4976 17674
rect 4754 16093 4788 17767
rect 5036 16093 5070 17860
rect 5224 16093 5258 17953
rect 4848 16093 4882 18046
rect 4660 16093 4694 18139
rect 6860 16093 6894 18232
rect 6672 16093 6706 18325
rect 6484 16093 6518 18418
rect 6296 16093 6330 18511
rect 6202 16093 6236 18604
rect 6108 16093 6142 18697
rect 6014 16093 6048 18790
rect 5920 16093 5954 18883
rect 4824 -826 4858 281
rect 6696 -826 6730 281
rect -1315 24166 -361 24200
rect 1115 24386 1283 24420
rect 1283 24102 2159 24136
rect 2125 24102 2159 24200
rect 1283 24102 1317 24420
rect 3635 24386 3803 24420
rect 3803 24102 4679 24136
rect 4645 24102 4679 24200
rect 3803 24102 3837 24420
rect 6155 24386 6323 24420
rect 6323 24102 7199 24136
rect 7165 24102 7199 24200
rect 6323 24102 6357 24420
rect 8675 24386 8843 24420
rect 8843 24102 9719 24136
rect 9685 24102 9719 24200
rect 8843 24102 8877 24420
rect 10915 23726 11033 23760
rect 9989 23506 10915 23540
rect 10915 23506 10949 23760
rect -883 2493 34 2527
rect -883 4193 34 4227
rect -883 5893 34 5927
rect -883 7593 34 7627
rect -883 9293 34 9327
rect -883 10993 34 11027
rect -883 12693 34 12727
rect -883 14393 34 14427
rect 11520 2493 12437 2527
rect 11520 4193 12437 4227
rect 11520 5893 12437 5927
rect 11520 7593 12437 7627
rect 11520 9293 12437 9327
rect 11520 10993 12437 11027
rect 11520 12693 12437 12727
rect 11520 14393 12437 14427
<< locali >>
rect 12345 -360 12437 24983
rect -883 -360 12437 -268
rect -883 24891 12437 24983
rect -883 -360 -791 24983
rect 12345 -360 12437 24983
rect 12705 -720 12797 25343
rect -1243 -720 12797 -628
rect -1243 25251 12797 25343
rect -1243 -720 -1151 25343
rect 12705 -720 12797 25343
rect -1243 25611 12797 25703
rect -1243 25611 12797 25703
rect 12869 -826 12903 25703
rect -1243 -826 12903 -792
rect 12869 -826 12903 25703
rect -1349 -932 12903 -898
rect -1349 -932 -1315 25703
rect 9935 23506 10043 23540
rect -361 22934 -253 22968
rect 467 20910 575 20944
rect 5291 1259 5399 1293
rect 5291 555 5399 589
use SUNSAR_SARBSSW_CV XB1 
transform -1 0 5777 0 1 0
box 5777 0 11501 2400
use SUNSAR_SARBSSW_CV XB2 
transform 1 0 5777 0 1 0
box 5777 0 11501 2400
use SUNSAR_CDAC8_CV XDAC1 
transform -1 0 5702 0 1 2493
box 5702 2493 11336 16127
use SUNSAR_CDAC8_CV XDAC2 
transform 1 0 5852 0 1 2493
box 5852 2493 11486 16127
use SUNSAR_SARDIGEX4_CV XA0 
transform 1 0 -523 0 1 19255
box -523 19255 737 24623
use SUNSAR_SARDIGEX4_CV XA1 
transform -1 0 1997 0 1 19255
box 1997 19255 3257 24623
use SUNSAR_SARDIGEX4_CV XA2 
transform 1 0 1997 0 1 19255
box 1997 19255 3257 24623
use SUNSAR_SARDIGEX4_CV XA3 
transform -1 0 4517 0 1 19255
box 4517 19255 5777 24623
use SUNSAR_SARDIGEX4_CV XA4 
transform 1 0 4517 0 1 19255
box 4517 19255 5777 24623
use SUNSAR_SARDIGEX4_CV XA5 
transform -1 0 7037 0 1 19255
box 7037 19255 8297 24623
use SUNSAR_SARDIGEX4_CV XA6 
transform 1 0 7037 0 1 19255
box 7037 19255 8297 24623
use SUNSAR_SARDIGEX4_CV XA7 
transform -1 0 9557 0 1 19255
box 9557 19255 10817 24623
use SUNSAR_SARDIGEX4_CV XA8 
transform 1 0 9557 0 1 19255
box 9557 19255 10817 24623
use SUNSAR_SARCMPX1_CV XA20 
transform -1 0 12077 0 1 19255
box 12077 19255 13337 24183
use SUNSAR_cut_M3M4_1x2 xcut0 
transform 1 0 7230 0 1 16127
box 7230 16127 7264 16219
use SUNSAR_cut_M3M4_2x1 xcut1 
transform 1 0 7230 0 1 16372
box 7230 16372 7322 16406
use SUNSAR_cut_M3M4_1x2 xcut2 
transform 1 0 4290 0 1 16127
box 4290 16127 4324 16219
use SUNSAR_cut_M3M4_2x1 xcut3 
transform 1 0 4290 0 1 16558
box 4290 16558 4382 16592
use SUNSAR_cut_M2M4_2x1 xcut4 
transform 1 0 11807 0 1 19942
box 11807 19942 11899 19976
use SUNSAR_cut_M4M5_2x1 xcut5 
transform 1 0 11807 0 1 16558
box 11807 16558 11903 16592
use SUNSAR_cut_M4M5_1x2 xcut6 
transform 1 0 11807 0 1 16728
box 11807 16728 11841 16824
use SUNSAR_cut_M3M4_2x1 xcut7 
transform 1 0 11887 0 1 22230
box 11887 22230 11979 22264
use SUNSAR_cut_M2M3_2x1 xcut8 
transform 1 0 11807 0 1 22230
box 11807 22230 11899 22264
use SUNSAR_cut_M4M5_2x1 xcut9 
transform 1 0 11945 0 1 16372
box 11945 16372 12041 16406
use SUNSAR_cut_M4M5_1x2 xcut10 
transform 1 0 11945 0 1 16728
box 11945 16728 11979 16824
use SUNSAR_cut_M3M4_1x2 xcut11 
transform 1 0 -345 0 1 16715
box -345 16715 -311 16807
use SUNSAR_cut_M2M3_1x2 xcut12 
transform 1 0 6954 0 1 16715
box 6954 16715 6988 16807
use SUNSAR_cut_M3M4_1x2 xcut13 
transform 1 0 4247 0 1 16808
box 4247 16808 4281 16900
use SUNSAR_cut_M2M3_1x2 xcut14 
transform 1 0 6390 0 1 16808
box 6390 16808 6424 16900
use SUNSAR_cut_M3M4_1x2 xcut15 
transform 1 0 2175 0 1 16901
box 2175 16901 2209 16993
use SUNSAR_cut_M2M3_1x2 xcut16 
transform 1 0 6578 0 1 16901
box 6578 16901 6612 16993
use SUNSAR_cut_M3M4_1x2 xcut17 
transform 1 0 1727 0 1 16994
box 1727 16994 1761 17086
use SUNSAR_cut_M2M3_1x2 xcut18 
transform 1 0 6766 0 1 16994
box 6766 16994 6800 17086
use SUNSAR_cut_M3M4_1x2 xcut19 
transform 1 0 0 0 1 17087
box 0 17087 34 17179
use SUNSAR_cut_M2M3_1x2 xcut20 
transform 1 0 4566 0 1 17087
box 4566 17087 4600 17179
use SUNSAR_cut_M3M4_1x2 xcut21 
transform 1 0 3959 0 1 17180
box 3959 17180 3993 17272
use SUNSAR_cut_M2M3_1x2 xcut22 
transform 1 0 5130 0 1 17180
box 5130 17180 5164 17272
use SUNSAR_cut_M3M4_1x2 xcut23 
transform 1 0 5040 0 1 17273
box 5040 17273 5074 17365
use SUNSAR_cut_M2M3_1x2 xcut24 
transform 1 0 5318 0 1 17273
box 5318 17273 5352 17365
use SUNSAR_cut_M3M4_1x2 xcut25 
transform 1 0 6479 0 1 17366
box 6479 17366 6513 17458
use SUNSAR_cut_M2M3_1x2 xcut26 
transform 1 0 5412 0 1 17366
box 5412 17366 5446 17458
use SUNSAR_cut_M3M4_1x2 xcut27 
transform 1 0 7560 0 1 17459
box 7560 17459 7594 17551
use SUNSAR_cut_M2M3_1x2 xcut28 
transform 1 0 5506 0 1 17459
box 5506 17459 5540 17551
use SUNSAR_cut_M3M4_1x2 xcut29 
transform 1 0 8999 0 1 17552
box 8999 17552 9033 17644
use SUNSAR_cut_M2M3_1x2 xcut30 
transform 1 0 5600 0 1 17552
box 5600 17552 5634 17644
use SUNSAR_cut_M3M4_1x2 xcut31 
transform 1 0 2520 0 1 17645
box 2520 17645 2554 17737
use SUNSAR_cut_M2M3_1x2 xcut32 
transform 1 0 4942 0 1 17645
box 4942 17645 4976 17737
use SUNSAR_cut_M3M4_1x2 xcut33 
transform 1 0 1439 0 1 17738
box 1439 17738 1473 17830
use SUNSAR_cut_M2M3_1x2 xcut34 
transform 1 0 4754 0 1 17738
box 4754 17738 4788 17830
use SUNSAR_cut_M3M4_1x2 xcut35 
transform 1 0 2591 0 1 17831
box 2591 17831 2625 17923
use SUNSAR_cut_M2M3_1x2 xcut36 
transform 1 0 5036 0 1 17831
box 5036 17831 5070 17923
use SUNSAR_cut_M3M4_1x2 xcut37 
transform 1 0 3888 0 1 17924
box 3888 17924 3922 18016
use SUNSAR_cut_M2M3_1x2 xcut38 
transform 1 0 5224 0 1 17924
box 5224 17924 5258 18016
use SUNSAR_cut_M3M4_1x2 xcut39 
transform 1 0 1368 0 1 18017
box 1368 18017 1402 18109
use SUNSAR_cut_M2M3_1x2 xcut40 
transform 1 0 4848 0 1 18017
box 4848 18017 4882 18109
use SUNSAR_cut_M3M4_1x2 xcut41 
transform 1 0 71 0 1 18110
box 71 18110 105 18202
use SUNSAR_cut_M2M3_1x2 xcut42 
transform 1 0 4660 0 1 18110
box 4660 18110 4694 18202
use SUNSAR_cut_M3M4_1x2 xcut43 
transform 1 0 150 0 1 18203
box 150 18203 184 18295
use SUNSAR_cut_M2M3_1x2 xcut44 
transform 1 0 6860 0 1 18203
box 6860 18203 6894 18295
use SUNSAR_cut_M3M4_1x2 xcut45 
transform 1 0 1290 0 1 18296
box 1290 18296 1324 18388
use SUNSAR_cut_M2M3_1x2 xcut46 
transform 1 0 6672 0 1 18296
box 6672 18296 6706 18388
use SUNSAR_cut_M3M4_1x2 xcut47 
transform 1 0 2670 0 1 18389
box 2670 18389 2704 18481
use SUNSAR_cut_M2M3_1x2 xcut48 
transform 1 0 6484 0 1 18389
box 6484 18389 6518 18481
use SUNSAR_cut_M3M4_1x2 xcut49 
transform 1 0 3810 0 1 18482
box 3810 18482 3844 18574
use SUNSAR_cut_M2M3_1x2 xcut50 
transform 1 0 6296 0 1 18482
box 6296 18482 6330 18574
use SUNSAR_cut_M3M4_1x2 xcut51 
transform 1 0 5190 0 1 18575
box 5190 18575 5224 18667
use SUNSAR_cut_M2M3_1x2 xcut52 
transform 1 0 6202 0 1 18575
box 6202 18575 6236 18667
use SUNSAR_cut_M3M4_1x2 xcut53 
transform 1 0 6330 0 1 18668
box 6330 18668 6364 18760
use SUNSAR_cut_M2M3_1x2 xcut54 
transform 1 0 6108 0 1 18668
box 6108 18668 6142 18760
use SUNSAR_cut_M3M4_1x2 xcut55 
transform 1 0 7710 0 1 18761
box 7710 18761 7744 18853
use SUNSAR_cut_M2M3_1x2 xcut56 
transform 1 0 6014 0 1 18761
box 6014 18761 6048 18853
use SUNSAR_cut_M3M4_1x2 xcut57 
transform 1 0 8850 0 1 18854
box 8850 18854 8884 18946
use SUNSAR_cut_M2M3_1x2 xcut58 
transform 1 0 5920 0 1 18854
box 5920 18854 5954 18946
use SUNSAR_cut_M1M4_2x2 xcut59 
transform 1 0 -145 0 1 24891
box -145 24891 -53 24983
use SUNSAR_cut_M1M4_2x2 xcut60 
transform 1 0 1527 0 1 24891
box 1527 24891 1619 24983
use SUNSAR_cut_M1M4_2x2 xcut61 
transform 1 0 2375 0 1 24891
box 2375 24891 2467 24983
use SUNSAR_cut_M1M4_2x2 xcut62 
transform 1 0 4047 0 1 24891
box 4047 24891 4139 24983
use SUNSAR_cut_M1M4_2x2 xcut63 
transform 1 0 4895 0 1 24891
box 4895 24891 4987 24983
use SUNSAR_cut_M1M4_2x2 xcut64 
transform 1 0 6567 0 1 24891
box 6567 24891 6659 24983
use SUNSAR_cut_M1M4_2x2 xcut65 
transform 1 0 7415 0 1 24891
box 7415 24891 7507 24983
use SUNSAR_cut_M1M4_2x2 xcut66 
transform 1 0 9087 0 1 24891
box 9087 24891 9179 24983
use SUNSAR_cut_M1M4_2x2 xcut67 
transform 1 0 9935 0 1 24891
box 9935 24891 10027 24983
use SUNSAR_cut_M1M4_2x2 xcut68 
transform 1 0 11607 0 1 24891
box 11607 24891 11699 24983
use SUNSAR_cut_M1M4_2x2 xcut69 
transform 1 0 4587 0 1 -360
box 4587 -360 4679 -268
use SUNSAR_cut_M1M4_2x2 xcut70 
transform 1 0 6875 0 1 -360
box 6875 -360 6967 -268
use SUNSAR_cut_M1M4_2x2 xcut71 
transform 1 0 251 0 1 25251
box 251 25251 343 25343
use SUNSAR_cut_M1M4_2x2 xcut72 
transform 1 0 1131 0 1 25251
box 1131 25251 1223 25343
use SUNSAR_cut_M1M4_2x2 xcut73 
transform 1 0 2771 0 1 25251
box 2771 25251 2863 25343
use SUNSAR_cut_M1M4_2x2 xcut74 
transform 1 0 3651 0 1 25251
box 3651 25251 3743 25343
use SUNSAR_cut_M1M4_2x2 xcut75 
transform 1 0 5291 0 1 25251
box 5291 25251 5383 25343
use SUNSAR_cut_M1M4_2x2 xcut76 
transform 1 0 6171 0 1 25251
box 6171 25251 6263 25343
use SUNSAR_cut_M1M4_2x2 xcut77 
transform 1 0 7811 0 1 25251
box 7811 25251 7903 25343
use SUNSAR_cut_M1M4_2x2 xcut78 
transform 1 0 8691 0 1 25251
box 8691 25251 8783 25343
use SUNSAR_cut_M1M4_2x2 xcut79 
transform 1 0 10331 0 1 25251
box 10331 25251 10423 25343
use SUNSAR_cut_M1M4_2x2 xcut80 
transform 1 0 11211 0 1 25251
box 11211 25251 11303 25343
use SUNSAR_cut_M1M4_2x2 xcut81 
transform 1 0 4191 0 1 -720
box 4191 -720 4283 -628
use SUNSAR_cut_M1M4_2x2 xcut82 
transform 1 0 7271 0 1 -720
box 7271 -720 7363 -628
use SUNSAR_cut_M1M4_2x2 xcut83 
transform 1 0 539 0 1 25611
box 539 25611 631 25703
use SUNSAR_cut_M1M4_2x2 xcut84 
transform 1 0 843 0 1 25611
box 843 25611 935 25703
use SUNSAR_cut_M1M4_2x2 xcut85 
transform 1 0 3059 0 1 25611
box 3059 25611 3151 25703
use SUNSAR_cut_M1M4_2x2 xcut86 
transform 1 0 3363 0 1 25611
box 3363 25611 3455 25703
use SUNSAR_cut_M1M4_2x2 xcut87 
transform 1 0 5579 0 1 25611
box 5579 25611 5671 25703
use SUNSAR_cut_M1M4_2x2 xcut88 
transform 1 0 5883 0 1 25611
box 5883 25611 5975 25703
use SUNSAR_cut_M1M4_2x2 xcut89 
transform 1 0 8099 0 1 25611
box 8099 25611 8191 25703
use SUNSAR_cut_M1M4_2x2 xcut90 
transform 1 0 8403 0 1 25611
box 8403 25611 8495 25703
use SUNSAR_cut_M1M4_2x2 xcut91 
transform 1 0 10619 0 1 25611
box 10619 25611 10711 25703
use SUNSAR_cut_M1M2_2x1 xcut92 
transform 1 0 4795 0 1 247
box 4795 247 4887 281
use SUNSAR_cut_M1M2_2x1 xcut93 
transform 1 0 4795 0 1 -826
box 4795 -826 4887 -792
use SUNSAR_cut_M1M2_2x1 xcut94 
transform 1 0 6667 0 1 247
box 6667 247 6759 281
use SUNSAR_cut_M1M2_2x1 xcut95 
transform 1 0 6667 0 1 -826
box 6667 -826 6759 -792
use SUNSAR_cut_M1M2_2x1 xcut96 
transform 1 0 -361 0 1 24166
box -361 24166 -269 24200
use SUNSAR_cut_M1M2_1x2 xcut97 
transform 1 0 -1349 0 1 24137
box -1349 24137 -1315 24229
use SUNSAR_cut_M1M4_2x1 xcut98 
transform 1 0 4847 0 1 -932
box 4847 -932 4939 -898
use SUNSAR_cut_M1M4_2x1 xcut99 
transform 1 0 6615 0 1 -932
box 6615 -932 6707 -898
use SUNSAR_cut_M1M3_2x1 xcut100 
transform 1 0 251 0 1 24403
box 251 24403 343 24437
use SUNSAR_cut_M1M3_2x1 xcut101 
transform 1 0 1727 0 1 24166
box 1727 24166 1819 24200
use SUNSAR_cut_M1M3_2x1 xcut102 
transform 1 0 2771 0 1 24403
box 2771 24403 2863 24437
use SUNSAR_cut_M1M3_2x1 xcut103 
transform 1 0 4247 0 1 24166
box 4247 24166 4339 24200
use SUNSAR_cut_M1M3_2x1 xcut104 
transform 1 0 5291 0 1 24403
box 5291 24403 5383 24437
use SUNSAR_cut_M1M3_2x1 xcut105 
transform 1 0 6767 0 1 24166
box 6767 24166 6859 24200
use SUNSAR_cut_M1M3_2x1 xcut106 
transform 1 0 7811 0 1 24403
box 7811 24403 7903 24437
use SUNSAR_cut_M1M3_2x1 xcut107 
transform 1 0 9287 0 1 24166
box 9287 24166 9379 24200
use SUNSAR_cut_M1M3_2x1 xcut108 
transform 1 0 -361 0 1 22934
box -361 22934 -269 22968
use SUNSAR_cut_M1M3_2x1 xcut109 
transform 1 0 1727 0 1 22934
box 1727 22934 1819 22968
use SUNSAR_cut_M1M3_2x1 xcut110 
transform 1 0 2159 0 1 22934
box 2159 22934 2251 22968
use SUNSAR_cut_M1M3_2x1 xcut111 
transform 1 0 4247 0 1 22934
box 4247 22934 4339 22968
use SUNSAR_cut_M1M3_2x1 xcut112 
transform 1 0 4679 0 1 22934
box 4679 22934 4771 22968
use SUNSAR_cut_M1M3_2x1 xcut113 
transform 1 0 6767 0 1 22934
box 6767 22934 6859 22968
use SUNSAR_cut_M1M3_2x1 xcut114 
transform 1 0 7199 0 1 22934
box 7199 22934 7291 22968
use SUNSAR_cut_M1M3_2x1 xcut115 
transform 1 0 9287 0 1 22934
box 9287 22934 9379 22968
use SUNSAR_cut_M1M3_2x1 xcut116 
transform 1 0 9719 0 1 22934
box 9719 22934 9811 22968
use SUNSAR_cut_M1M2_2x1 xcut117 
transform 1 0 1115 0 1 24386
box 1115 24386 1207 24420
use SUNSAR_cut_M1M2_2x1 xcut118 
transform 1 0 2159 0 1 24166
box 2159 24166 2251 24200
use SUNSAR_cut_M1M2_2x1 xcut119 
transform 1 0 3635 0 1 24386
box 3635 24386 3727 24420
use SUNSAR_cut_M1M2_2x1 xcut120 
transform 1 0 4679 0 1 24166
box 4679 24166 4771 24200
use SUNSAR_cut_M1M2_2x1 xcut121 
transform 1 0 6155 0 1 24386
box 6155 24386 6247 24420
use SUNSAR_cut_M1M2_2x1 xcut122 
transform 1 0 7199 0 1 24166
box 7199 24166 7291 24200
use SUNSAR_cut_M1M2_2x1 xcut123 
transform 1 0 8675 0 1 24386
box 8675 24386 8767 24420
use SUNSAR_cut_M1M2_2x1 xcut124 
transform 1 0 9719 0 1 24166
box 9719 24166 9811 24200
use SUNSAR_cut_M1M3_2x1 xcut125 
transform 1 0 -361 0 1 20734
box -361 20734 -269 20768
use SUNSAR_cut_M1M3_2x1 xcut126 
transform 1 0 1727 0 1 20734
box 1727 20734 1819 20768
use SUNSAR_cut_M1M3_2x1 xcut127 
transform 1 0 2159 0 1 20734
box 2159 20734 2251 20768
use SUNSAR_cut_M1M3_2x1 xcut128 
transform 1 0 4247 0 1 20734
box 4247 20734 4339 20768
use SUNSAR_cut_M1M3_2x1 xcut129 
transform 1 0 4679 0 1 20734
box 4679 20734 4771 20768
use SUNSAR_cut_M1M3_2x1 xcut130 
transform 1 0 6767 0 1 20734
box 6767 20734 6859 20768
use SUNSAR_cut_M1M3_2x1 xcut131 
transform 1 0 7199 0 1 20734
box 7199 20734 7291 20768
use SUNSAR_cut_M1M3_2x1 xcut132 
transform 1 0 9287 0 1 20734
box 9287 20734 9379 20768
use SUNSAR_cut_M1M3_2x1 xcut133 
transform 1 0 9719 0 1 20734
box 9719 20734 9811 20768
use SUNSAR_cut_M1M3_2x1 xcut134 
transform 1 0 467 0 1 20910
box 467 20910 559 20944
use SUNSAR_cut_M1M3_2x1 xcut135 
transform 1 0 899 0 1 20910
box 899 20910 991 20944
use SUNSAR_cut_M1M3_2x1 xcut136 
transform 1 0 2987 0 1 20910
box 2987 20910 3079 20944
use SUNSAR_cut_M1M3_2x1 xcut137 
transform 1 0 3419 0 1 20910
box 3419 20910 3511 20944
use SUNSAR_cut_M1M3_2x1 xcut138 
transform 1 0 5507 0 1 20910
box 5507 20910 5599 20944
use SUNSAR_cut_M1M3_2x1 xcut139 
transform 1 0 5939 0 1 20910
box 5939 20910 6031 20944
use SUNSAR_cut_M1M3_2x1 xcut140 
transform 1 0 8027 0 1 20910
box 8027 20910 8119 20944
use SUNSAR_cut_M1M3_2x1 xcut141 
transform 1 0 8459 0 1 20910
box 8459 20910 8551 20944
use SUNSAR_cut_M1M3_2x1 xcut142 
transform 1 0 10547 0 1 20910
box 10547 20910 10639 20944
use SUNSAR_cut_M1M3_2x1 xcut143 
transform 1 0 11607 0 1 20971
box 11607 20971 11699 21005
use SUNSAR_cut_M1M3_2x1 xcut144 
transform 1 0 11211 0 1 21411
box 11211 21411 11303 21445
use SUNSAR_cut_M1M3_2x1 xcut145 
transform 1 0 10979 0 1 23638
box 10979 23638 11071 23672
use SUNSAR_cut_M1M3_2x1 xcut146 
transform 1 0 9719 0 1 23110
box 9719 23110 9811 23144
use SUNSAR_cut_M1M3_2x1 xcut147 
transform 1 0 10995 0 1 23902
box 10995 23902 11087 23936
use SUNSAR_cut_M1M3_2x1 xcut148 
transform 1 0 10347 0 1 24403
box 10347 24403 10439 24437
use SUNSAR_cut_M1M2_2x1 xcut149 
transform 1 0 10995 0 1 23726
box 10995 23726 11087 23760
use SUNSAR_cut_M1M2_2x1 xcut150 
transform 1 0 9951 0 1 23506
box 9951 23506 10043 23540
use SUNSAR_cut_M4M5_1x2 xcut151 
transform 1 0 5227 0 1 555
box 5227 555 5261 651
use SUNSAR_cut_M4M5_1x2 xcut152 
transform 1 0 5227 0 1 2431
box 5227 2431 5261 2527
use SUNSAR_cut_M1M4_2x1 xcut153 
transform 1 0 6155 0 1 555
box 6155 555 6247 589
use SUNSAR_cut_M4M5_1x2 xcut154 
transform 1 0 6293 0 1 555
box 6293 555 6327 651
use SUNSAR_cut_M4M5_1x2 xcut155 
transform 1 0 6293 0 1 2431
box 6293 2431 6327 2527
use SUNSAR_cut_M1M3_2x1 xcut156 
transform 1 0 5291 0 1 1259
box 5291 1259 5383 1293
use SUNSAR_cut_M1M3_2x1 xcut157 
transform 1 0 6155 0 1 555
box 6155 555 6247 589
use SUNSAR_cut_M1M4_2x1 xcut158 
transform 1 0 5291 0 1 555
box 5291 555 5383 589
use SUNSAR_cut_M1M4_2x1 xcut159 
transform 1 0 6155 0 1 1259
box 6155 1259 6247 1293
use SUNSAR_cut_M1M3_2x1 xcut160 
transform 1 0 -361 0 1 20910
box -361 20910 -269 20944
use SUNSAR_cut_M1M2_2x2 xcut161 
transform 1 0 -883 0 1 2527
box -883 2527 -791 2619
use SUNSAR_cut_M1M2_2x2 xcut162 
transform 1 0 -883 0 1 4227
box -883 4227 -791 4319
use SUNSAR_cut_M1M2_2x2 xcut163 
transform 1 0 -883 0 1 5927
box -883 5927 -791 6019
use SUNSAR_cut_M1M2_2x2 xcut164 
transform 1 0 -883 0 1 7627
box -883 7627 -791 7719
use SUNSAR_cut_M1M2_2x2 xcut165 
transform 1 0 -883 0 1 9327
box -883 9327 -791 9419
use SUNSAR_cut_M1M2_2x2 xcut166 
transform 1 0 -883 0 1 11027
box -883 11027 -791 11119
use SUNSAR_cut_M1M2_2x2 xcut167 
transform 1 0 -883 0 1 12727
box -883 12727 -791 12819
use SUNSAR_cut_M1M2_2x2 xcut168 
transform 1 0 -883 0 1 14427
box -883 14427 -791 14519
use SUNSAR_cut_M1M2_1x2 xcut169 
transform 1 0 12403 0 1 2493
box 12403 2493 12437 2585
use SUNSAR_cut_M1M2_1x2 xcut170 
transform 1 0 12403 0 1 4193
box 12403 4193 12437 4285
use SUNSAR_cut_M1M2_1x2 xcut171 
transform 1 0 12403 0 1 5893
box 12403 5893 12437 5985
use SUNSAR_cut_M1M2_1x2 xcut172 
transform 1 0 12403 0 1 7593
box 12403 7593 12437 7685
use SUNSAR_cut_M1M2_1x2 xcut173 
transform 1 0 12403 0 1 9293
box 12403 9293 12437 9385
use SUNSAR_cut_M1M2_1x2 xcut174 
transform 1 0 12403 0 1 10993
box 12403 10993 12437 11085
use SUNSAR_cut_M1M2_1x2 xcut175 
transform 1 0 12403 0 1 12693
box 12403 12693 12437 12785
use SUNSAR_cut_M1M2_1x2 xcut176 
transform 1 0 12403 0 1 14393
box 12403 14393 12437 14485
<< labels >>
flabel m3 s -345 16778 -311 21526 0 FreeSans 400 0 0 0 D<8>
port 6 nsew signal bidirectional
flabel m3 s 3959 17243 3993 21541 0 FreeSans 400 0 0 0 D<5>
port 9 nsew signal bidirectional
flabel m3 s 5040 17336 5074 21541 0 FreeSans 400 0 0 0 D<4>
port 10 nsew signal bidirectional
flabel m3 s 6479 17429 6513 21541 0 FreeSans 400 0 0 0 D<3>
port 11 nsew signal bidirectional
flabel m3 s 7560 17522 7594 21541 0 FreeSans 400 0 0 0 D<2>
port 12 nsew signal bidirectional
flabel m3 s 8999 17615 9033 21541 0 FreeSans 400 0 0 0 D<1>
port 13 nsew signal bidirectional
flabel m3 s 2520 17708 2554 21541 0 FreeSans 400 0 0 0 D<6>
port 8 nsew signal bidirectional
flabel m3 s 1439 17801 1473 21541 0 FreeSans 400 0 0 0 D<7>
port 7 nsew signal bidirectional
flabel locali s 12345 -360 12437 24983 0 FreeSans 400 0 0 0 AVSS
port 20 nsew signal bidirectional
flabel locali s 12705 -720 12797 25343 0 FreeSans 400 0 0 0 AVDD
port 19 nsew signal bidirectional
flabel locali s -1243 25611 12797 25703 0 FreeSans 400 0 0 0 VREF
port 18 nsew signal bidirectional
flabel locali s 12869 -826 12903 25703 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew signal bidirectional
flabel locali s 9935 23506 10043 23540 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel m3 s 5291 115 5383 149 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel m3 s 6171 115 6263 149 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s -361 22934 -253 22968 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew signal bidirectional
flabel locali s 467 20910 575 20944 0 FreeSans 400 0 0 0 EN
port 15 nsew signal bidirectional
flabel locali s 5291 1259 5399 1293 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 5291 555 5399 589 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel m3 s 10080 21541 10114 21633 0 FreeSans 400 0 0 0 D<0>
port 14 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -1349 -932 12903 25703
<< end >>
