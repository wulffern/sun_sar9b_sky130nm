magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 1260 352
<< locali >>
rect 415 115 449 149
rect 415 203 449 237
rect 811 203 845 237
rect 432 291 516 325
rect 516 291 828 325
rect 516 291 550 325
rect 710 27 828 61
rect 710 203 828 237
rect 710 27 744 237
rect 378 203 882 237
rect 162 159 270 193
rect 990 247 1098 281
rect 162 247 270 281
rect 162 71 270 105
rect 378 291 486 325
rect 1206 154 1314 198
rect -54 154 54 198
<< poly >>
rect 162 167 1098 185
rect 162 79 1098 97
<< m3 >>
rect 774 0 874 352
rect 378 0 478 352
rect 774 0 874 352
rect 378 0 478 352
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 88
box 0 88 630 264
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 176
box 0 176 630 352
use SUNSAR_PCHDL MP2 
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNSAR_PCHDL MP0 
transform 1 0 630 0 1 88
box 630 88 1260 264
use SUNSAR_PCHDL MP1 
transform 1 0 630 0 1 176
box 630 176 1260 352
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 115
box 774 115 874 153
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 115
box 774 115 874 153
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 27
box 378 27 478 65
<< labels >>
flabel locali s 162 159 270 193 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 990 247 1098 281 0 FreeSans 400 0 0 0 CN
port 3 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 400 0 0 0 C
port 2 nsew signal bidirectional
flabel locali s 162 71 270 105 0 FreeSans 400 0 0 0 RN
port 4 nsew signal bidirectional
flabel locali s 378 291 486 325 0 FreeSans 400 0 0 0 Y
port 5 nsew signal bidirectional
flabel locali s 1206 154 1314 198 0 FreeSans 400 0 0 0 BULKP
port 6 nsew signal bidirectional
flabel locali s -54 154 54 198 0 FreeSans 400 0 0 0 BULKN
port 7 nsew signal bidirectional
flabel m3 s 774 0 874 352 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 378 0 478 352 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 352
<< end >>
