magic
tech sky130A
timestamp 1712959200
<< checkpaint >>
rect 0 0 92 92
<< metal1 >>
rect 0 86 92 92
rect 0 58 6 86
rect 34 58 58 86
rect 86 58 92 86
rect 0 34 92 58
rect 0 6 6 34
rect 34 6 58 34
rect 86 6 92 34
rect 0 0 92 6
<< via1 >>
rect 6 58 34 86
rect 58 58 86 86
rect 6 6 34 34
rect 58 6 86 34
<< metal2 >>
rect 0 86 92 92
rect 0 58 6 86
rect 34 58 58 86
rect 86 58 92 86
rect 0 34 92 58
rect 0 6 6 34
rect 34 6 58 34
rect 86 6 92 34
rect 0 0 92 6
<< via2 >>
rect 6 58 34 86
rect 58 58 86 86
rect 6 6 34 34
rect 58 6 86 34
<< metal3 >>
rect 0 86 92 92
rect 0 58 6 86
rect 34 58 58 86
rect 86 58 92 86
rect 0 34 92 58
rect 0 6 6 34
rect 34 6 58 34
rect 86 6 92 34
rect 0 0 92 6
<< properties >>
string FIXED_BBOX 0 0 92 92
<< end >>
