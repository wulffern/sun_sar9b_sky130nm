magic
tech sky130B
magscale 1 2
timestamp 1708642800
<< checkpaint >>
rect 0 0 2520 3872
<< locali >>
rect 1656 582 1824 650
rect 1824 778 2040 846
rect 1824 582 1892 846
rect 1980 846 2088 914
rect 1656 934 1824 1002
rect 1824 1374 2088 1442
rect 1824 3310 2088 3378
rect 1824 934 1892 3378
rect 432 1902 600 1970
rect 600 934 864 1002
rect 600 934 668 1970
rect 480 2714 600 2782
rect 600 934 864 1002
rect 600 934 668 2782
rect 432 2782 540 2850
rect 864 1462 1032 1530
rect 864 1990 1032 2058
rect 1032 1462 1100 2058
rect 864 2870 1032 2938
rect 864 3398 1032 3466
rect 1032 2870 1100 3466
rect 432 3662 600 3730
rect 600 3398 864 3466
rect 600 3398 668 3730
rect 324 1198 540 1266
rect 324 494 540 562
rect 756 3750 972 3818
rect 756 3398 972 3466
<< m1 >>
rect 2088 1902 2256 1970
rect 2088 2782 2256 2850
rect 1656 582 2256 650
rect 2256 582 2324 2850
rect 480 1306 600 1374
rect 600 582 864 650
rect 600 582 668 1374
rect 432 1374 540 1442
rect 432 3310 600 3378
rect 600 2782 2088 2850
rect 600 2782 668 3378
rect 432 2254 600 2322
rect 600 1990 864 2058
rect 600 1990 668 2322
rect 1656 2342 1824 2410
rect 1824 1726 2088 1794
rect 1824 2606 2088 2674
rect 1824 1726 1892 2674
rect 1656 3750 1824 3818
rect 1824 3134 2088 3202
rect 1824 3134 1892 3818
<< m3 >>
rect 1548 0 1732 3872
rect 756 0 940 3872
rect 1548 0 1732 3872
rect 756 0 940 3872
use SUNSAR_TAPCELLB_CV XA0 
transform 1 0 0 0 1 0
box 0 0 2520 352
use SUNSAR_IVX1_CV XA1 
transform 1 0 0 0 1 352
box 0 352 2520 704
use SUNSAR_IVX1_CV XA2 
transform 1 0 0 0 1 704
box 0 704 2520 1056
use SUNSAR_IVTRIX1_CV XA3 
transform 1 0 0 0 1 1056
box 0 1056 2520 1584
use SUNSAR_IVTRIX1_CV XA4 
transform 1 0 0 0 1 1584
box 0 1584 2520 2112
use SUNSAR_IVX1_CV XA5 
transform 1 0 0 0 1 2112
box 0 2112 2520 2464
use SUNSAR_IVTRIX1_CV XA6 
transform 1 0 0 0 1 2464
box 0 2464 2520 2992
use SUNSAR_IVTRIX1_CV XA7 
transform 1 0 0 0 1 2992
box 0 2992 2520 3520
use SUNSAR_IVX1_CV XA8 
transform 1 0 0 0 1 3520
box 0 3520 2520 3872
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 1980 0 1 1902
box 1980 1902 2164 1970
use SUNSAR_cut_M1M2_2x1 xcut1 
transform 1 0 1980 0 1 2782
box 1980 2782 2164 2850
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 1548 0 1 582
box 1548 582 1732 650
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 324 0 1 1374
box 324 1374 508 1442
use SUNSAR_cut_M1M2_2x1 xcut4 
transform 1 0 756 0 1 582
box 756 582 940 650
use SUNSAR_cut_M1M2_2x1 xcut5 
transform 1 0 324 0 1 3310
box 324 3310 508 3378
use SUNSAR_cut_M1M2_2x1 xcut6 
transform 1 0 1980 0 1 2782
box 1980 2782 2164 2850
use SUNSAR_cut_M1M2_2x1 xcut7 
transform 1 0 324 0 1 2254
box 324 2254 508 2322
use SUNSAR_cut_M1M2_2x1 xcut8 
transform 1 0 756 0 1 1990
box 756 1990 940 2058
use SUNSAR_cut_M1M2_2x1 xcut9 
transform 1 0 1548 0 1 2342
box 1548 2342 1732 2410
use SUNSAR_cut_M1M2_2x1 xcut10 
transform 1 0 1980 0 1 1726
box 1980 1726 2164 1794
use SUNSAR_cut_M1M2_2x1 xcut11 
transform 1 0 1980 0 1 2606
box 1980 2606 2164 2674
use SUNSAR_cut_M1M2_2x1 xcut12 
transform 1 0 1548 0 1 3750
box 1548 3750 1732 3818
use SUNSAR_cut_M1M2_2x1 xcut13 
transform 1 0 1980 0 1 3134
box 1980 3134 2164 3202
<< labels >>
flabel locali s 324 1198 540 1266 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 324 494 540 562 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 756 3750 972 3818 0 FreeSans 400 0 0 0 Q
port 3 nsew signal bidirectional
flabel locali s 756 3398 972 3466 0 FreeSans 400 0 0 0 QN
port 4 nsew signal bidirectional
flabel m3 s 1548 0 1732 3872 0 FreeSans 400 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel m3 s 756 0 940 3872 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 3872
<< end >>
