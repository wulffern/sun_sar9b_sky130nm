magic
tech sky130A
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 136 68
<< locali >>
rect 0 0 68 68
rect 0 0 68 68
rect 68 0 204 68
rect 68 0 204 68
<< rlocali >>
rect 68 0 136 68
<< labels >>
flabel locali s 0 0 68 68 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 68 0 204 68 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 136 68
<< end >>
