magic
tech sky130A
timestamp 1708968222
<< poly >>
rect 162 79 1098 97
<< locali >>
rect 378 115 486 149
rect 828 115 946 149
rect -54 66 54 110
rect 912 105 946 115
rect 912 71 1044 105
rect 1206 66 1314 110
<< metal3 >>
rect 378 0 470 176
rect 774 0 866 176
use SUNSAR_NCHDL  MN0
timestamp 1708902000
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNSAR_PCHDL  MP0
timestamp 1708902000
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNSAR_cut_M1M4_2x1  xcut0
timestamp 1708902000
transform 1 0 774 0 1 27
box 0 0 92 34
use SUNSAR_cut_M1M4_2x1  xcut1
timestamp 1708902000
transform 1 0 378 0 1 27
box 0 0 92 34
<< labels >>
flabel locali s 378 115 486 149 0 FreeSans 200 0 0 0 Y
port 1 nsew signal bidirectional
flabel locali s 1206 66 1314 110 0 FreeSans 200 0 0 0 BULKP
port 2 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 200 0 0 0 BULKN
port 3 nsew signal bidirectional
flabel metal3 s 774 0 866 176 0 FreeSans 200 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel metal3 s 378 0 470 176 0 FreeSans 200 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
