magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 68 34
<< locali >>
rect 0 0 34 34
rect 0 0 34 34
rect 34 0 102 34
rect 34 0 102 34
<< rlocali >>
rect 34 0 68 34
<< labels >>
flabel locali s 0 0 34 34 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 34 0 102 34 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 68 34
<< end >>
