magic
tech sky130A
magscale 1 2
timestamp 1708902000
<< checkpaint >>
rect 0 0 2520 880
<< locali >>
rect 432 670 600 738
rect 600 406 864 474
rect 600 406 668 738
rect 324 142 540 210
rect 324 318 540 386
rect 756 758 972 826
rect 2412 132 2628 220
rect -108 132 108 220
<< m3 >>
rect 1548 0 1732 880
rect 756 0 940 880
rect 1548 0 1732 880
rect 756 0 940 880
use SUNSAR_NDX1_CV XA1 
transform 1 0 0 0 1 0
box 0 0 2520 528
use SUNSAR_IVX1_CV XA2 
transform 1 0 0 0 1 528
box 0 528 2520 880
<< labels >>
flabel locali s 324 142 540 210 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 324 318 540 386 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 756 758 972 826 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 4 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 5 nsew signal bidirectional
flabel m3 s 1548 0 1732 880 0 FreeSans 400 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel m3 s 756 0 940 880 0 FreeSans 400 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 880
<< end >>
