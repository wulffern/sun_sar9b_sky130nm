magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 5724 2400
<< m1 >>
rect 1494 819 1710 853
rect 1548 291 1632 325
rect 1632 423 1764 457
rect 1632 291 1666 457
rect 216 1303 300 1337
rect 300 1435 1152 1469
rect 300 1303 334 1469
rect 936 863 1020 897
rect 1020 1100 1548 1134
rect 1020 863 1054 1134
rect 432 467 516 501
rect 516 643 1152 677
rect 516 467 550 677
<< locali >>
rect 0 1298 84 1332
rect 84 1562 720 1596
rect 84 1298 118 1596
rect 314 115 432 149
rect 314 291 432 325
rect 314 467 432 501
rect 314 643 432 677
rect 314 819 432 853
rect 314 995 432 1029
rect 314 1171 432 1205
rect 314 1347 432 1381
rect 314 115 348 1381
rect 199 71 233 633
rect 199 775 233 1337
rect 432 27 516 61
rect 432 203 516 237
rect 432 379 516 413
rect 432 555 516 589
rect 516 27 550 589
rect 432 731 516 765
rect 432 907 516 941
rect 432 1083 516 1117
rect 432 1259 516 1293
rect 516 731 550 1293
rect 882 247 990 281
rect 1710 423 1818 457
rect 378 555 486 589
rect 378 1259 486 1293
<< m2 >>
rect 936 775 1020 809
rect 1020 308 1152 342
rect 1020 308 1054 809
rect 716 907 1152 941
rect 216 423 716 457
rect 716 423 750 941
rect 1548 555 1632 589
rect 1632 -20 2192 14
rect 1632 -20 1666 589
<< m3 >>
rect 2078 1340 3924 1374
rect 1760 819 2078 853
rect 2078 819 2112 1374
rect 386 113 486 151
rect 806 1433 906 1471
rect 1494 0 1594 2400
rect 1098 0 1198 2400
rect 1494 0 1594 2400
rect 1098 0 1198 2400
use SUNSAR_NCHDLR M1 
transform 1 0 0 0 1 0
box 0 0 720 176
use SUNSAR_NCHDLR M2 
transform 1 0 0 0 1 176
box 0 176 720 352
use SUNSAR_NCHDLR M3 
transform 1 0 0 0 1 352
box 0 352 720 528
use SUNSAR_NCHDLR M4 
transform 1 0 0 0 1 528
box 0 528 720 704
use SUNSAR_NCHDLR M5 
transform 1 0 0 0 1 704
box 0 704 720 880
use SUNSAR_NCHDLR M6 
transform 1 0 0 0 1 880
box 0 880 720 1056
use SUNSAR_NCHDLR M7 
transform 1 0 0 0 1 1056
box 0 1056 720 1232
use SUNSAR_NCHDLR M8 
transform 1 0 0 0 1 1232
box 0 1232 720 1408
use SUNSAR_TAPCELLB_CV XA5b 
transform 1 0 720 0 1 0
box 720 0 1980 176
use SUNSAR_IVX1_CV XA0 
transform 1 0 720 0 1 176
box 720 176 1980 352
use SUNSAR_TGPD_CV XA3 
transform 1 0 720 0 1 352
box 720 352 1980 704
use SUNSAR_SARBSSWCTRL_CV XA4 
transform 1 0 720 0 1 704
box 720 704 1980 968
use SUNSAR_TIEH_CV XA1 
transform 1 0 720 0 1 968
box 720 968 1980 1144
use SUNSAR_TAPCELLB_CV XA7 
transform 1 0 720 0 1 1144
box 720 1144 1980 1320
use SUNSAR_TIEL_CV XA2 
transform 1 0 720 0 1 1320
box 720 1320 1980 1496
use SUNSAR_TAPCELLB_CV XA5 
transform 1 0 720 0 1 1496
box 720 1496 1980 1672
use SUNSAR_CAP_BSSW5_CV XCAPB1 
transform 1 0 2088 0 1 0
box 2088 0 5724 2400
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 1494 0 1 819
box 1494 819 1586 853
use SUNSAR_cut_M2M4_2x1 xcut1 
transform 1 0 1710 0 1 819
box 1710 819 1810 857
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 1494 0 1 291
box 1494 291 1586 325
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 1710 0 1 423
box 1710 423 1802 457
use SUNSAR_cut_M1M3_2x1 xcut4 
transform 1 0 882 0 1 775
box 882 775 974 809
use SUNSAR_cut_M1M3_2x1 xcut5 
transform 1 0 1098 0 1 308
box 1098 308 1190 342
use SUNSAR_cut_M1M2_2x1 xcut6 
transform 1 0 162 0 1 1303
box 162 1303 254 1337
use SUNSAR_cut_M1M2_2x1 xcut7 
transform 1 0 1098 0 1 1435
box 1098 1435 1190 1469
use SUNSAR_cut_M1M2_2x1 xcut8 
transform 1 0 882 0 1 863
box 882 863 974 897
use SUNSAR_cut_M1M2_2x1 xcut9 
transform 1 0 1494 0 1 1100
box 1494 1100 1586 1134
use SUNSAR_cut_M1M2_2x1 xcut10 
transform 1 0 378 0 1 467
box 378 467 470 501
use SUNSAR_cut_M1M2_2x1 xcut11 
transform 1 0 1098 0 1 643
box 1098 643 1190 677
use SUNSAR_cut_M1M3_2x1 xcut12 
transform 1 0 1114 0 1 907
box 1114 907 1206 941
use SUNSAR_cut_M1M3_2x1 xcut13 
transform 1 0 178 0 1 423
box 178 423 270 457
use SUNSAR_cut_M1M3_2x1 xcut14 
transform 1 0 1494 0 1 555
box 1494 555 1586 589
use SUNSAR_cut_M3M4_2x1 xcut15 
transform 1 0 2142 0 1 -20
box 2142 -20 2242 18
use SUNSAR_cut_M1M4_2x1 xcut16 
transform 1 0 386 0 1 113
box 386 113 486 151
use SUNSAR_cut_M2M4_2x1 xcut17 
transform 1 0 806 0 1 1433
box 806 1433 906 1471
<< labels >>
flabel m3 s 386 113 486 151 0 FreeSans 400 0 0 0 VI
port 1 nsew signal bidirectional
flabel m3 s 806 1433 906 1471 0 FreeSans 400 0 0 0 TIE_L
port 4 nsew signal bidirectional
flabel locali s 882 247 990 281 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 1710 423 1818 457 0 FreeSans 400 0 0 0 CKN
port 3 nsew signal bidirectional
flabel locali s 378 555 486 589 0 FreeSans 400 0 0 0 VO1
port 5 nsew signal bidirectional
flabel locali s 378 1259 486 1293 0 FreeSans 400 0 0 0 VO2
port 6 nsew signal bidirectional
flabel m3 s 1494 0 1594 2400 0 FreeSans 400 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel m3 s 1098 0 1198 2400 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 5724 2400
<< end >>
