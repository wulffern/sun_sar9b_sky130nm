magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 3636 2400
<< m3 >>
rect -10 380 1836 414
rect -10 860 1836 894
rect -10 1340 1836 1374
rect -10 1820 1836 1854
rect -10 2300 1836 2334
rect -10 380 24 2334
rect 1836 -20 3648 14
rect 1836 460 3648 494
rect 1836 940 3648 974
rect 1836 1420 3648 1454
rect 1836 1900 3648 1934
rect 3648 -20 3682 1934
rect 54 1340 3618 1380
rect 54 -20 3618 20
use SUNSAR_CAP_BSSW_CV XCAPB0 
transform 1 0 0 0 1 0
box 0 0 3636 480
use SUNSAR_CAP_BSSW_CV XCAPB1 
transform 1 0 0 0 1 480
box 0 480 3636 960
use SUNSAR_CAP_BSSW_CV XCAPB2 
transform 1 0 0 0 1 960
box 0 960 3636 1440
use SUNSAR_CAP_BSSW_CV XCAPB3 
transform 1 0 0 0 1 1440
box 0 1440 3636 1920
use SUNSAR_CAP_BSSW_CV XCAPB4 
transform 1 0 0 0 1 1920
box 0 1920 3636 2400
<< labels >>
flabel m3 s 54 1340 3618 1380 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel m3 s 54 -20 3618 20 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3636 2400
<< end >>
