magic
tech sky130B
magscale 1 2
timestamp 1681077600
<< checkpaint >>
rect 0 0 2520 2464
<< locali >>
rect 834 234 894 2230
rect 864 234 1032 294
rect 1032 58 1656 118
rect 1032 58 1092 294
rect 402 498 462 1966
rect 2058 498 2118 2318
rect 1626 234 1686 2406
rect 756 2346 1764 2406
rect 1656 2346 1824 2406
rect 1824 2258 2088 2318
rect 1824 2258 1884 2406
rect 834 234 894 470
rect 834 586 894 822
rect 834 938 894 1174
rect 834 1290 894 1526
rect 834 1642 894 1878
rect 834 1994 894 2230
rect 1626 234 1686 470
rect 1626 586 1686 822
rect 1626 938 1686 1174
rect 1626 1290 1686 1526
rect 1626 1642 1686 1878
rect 1626 1994 1686 2230
rect 2412 132 2628 220
rect -108 132 108 220
rect 324 2258 540 2318
rect 324 146 540 206
rect 324 498 540 558
<< poly >>
rect 324 158 2196 194
<< m3 >>
rect 1548 0 1748 2464
rect 756 0 956 2464
rect 1548 0 1748 2464
rect 756 0 956 2464
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNSAR_NCHDL MN2 
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNSAR_NCHDL MN3 
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNSAR_NCHDL MN4 
transform 1 0 0 0 1 1408
box 0 1408 1260 1760
use SUNSAR_NCHDL MN5 
transform 1 0 0 0 1 1760
box 0 1760 1260 2112
use SUNSAR_NCHDL MN6 
transform 1 0 0 0 1 2112
box 0 2112 1260 2464
use SUNSAR_PCHDL MP0 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1_DMY 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNSAR_PCHDL MP2_DMY 
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNSAR_PCHDL MP3_DMY 
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use SUNSAR_PCHDL MP4_DMY 
transform 1 0 1260 0 1 1408
box 1260 1408 2520 1760
use SUNSAR_PCHDL MP5_DMY 
transform 1 0 1260 0 1 1760
box 1260 1760 2520 2112
use SUNSAR_PCHDL MP6_DMY 
transform 1 0 1260 0 1 2112
box 1260 2112 2520 2464
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 234
box 1548 234 1748 310
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 756 0 1 58
box 756 58 956 134
<< labels >>
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 4 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 5 nsew signal bidirectional
flabel locali s 324 2258 540 2318 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 CKN
port 3 nsew signal bidirectional
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 CI
port 1 nsew signal bidirectional
flabel m3 s 1548 0 1748 2464 0 FreeSans 400 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel m3 s 756 0 956 2464 0 FreeSans 400 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 2464
<< end >>
