magic
tech sky130B
timestamp 1708692311
<< locali >>
rect 378 2051 486 2085
rect 216 2007 334 2041
rect 300 1909 334 2007
rect 300 1875 486 1909
rect 912 1831 1044 1865
rect 162 1655 270 1689
rect 216 1479 270 1513
rect 240 1445 334 1479
rect 300 1073 334 1445
rect 432 1083 550 1117
rect 216 1039 334 1073
rect 162 687 270 721
rect 300 589 334 1039
rect 516 853 550 1083
rect 432 819 550 853
rect 912 809 946 1831
rect 912 775 1044 809
rect 912 589 946 775
rect 300 555 432 589
rect 828 555 946 589
rect 990 511 1044 545
rect 912 477 1020 511
rect 912 325 946 477
rect 828 291 946 325
rect 162 247 270 281
<< metal1 >>
rect 828 2051 946 2085
rect 432 1875 550 1909
rect 216 1831 270 1865
rect 240 1797 334 1831
rect 98 1655 216 1689
rect 98 369 132 1655
rect 300 1479 334 1797
rect 516 1557 550 1875
rect 912 1777 946 2051
rect 912 1743 1044 1777
rect 432 1523 550 1557
rect 990 1479 1162 1513
rect 300 1445 1020 1479
rect 912 1391 1044 1425
rect 912 1293 946 1391
rect 828 1259 946 1293
rect 216 1215 334 1249
rect 300 1117 334 1215
rect 300 1083 432 1117
rect 912 985 946 1259
rect 1128 1073 1162 1479
rect 1044 1039 1162 1073
rect 912 951 1044 985
rect 216 775 270 809
rect 240 741 334 775
rect 300 413 334 741
rect 300 379 432 413
rect 98 335 216 369
rect 1128 325 1162 1039
rect 828 291 1162 325
<< metal3 >>
rect 378 0 470 2112
rect 774 0 866 2112
use SUNSAR_TAPCELLB_CV  XA0
timestamp 1708692311
transform 1 0 0 0 1 0
box -90 -66 1350 242
use SUNSAR_NDX1_CV  XA1
timestamp 1708692311
transform 1 0 0 0 1 176
box -90 -66 1350 330
use SUNSAR_IVX1_CV  XA2
timestamp 1708692311
transform 1 0 0 0 1 440
box -90 -66 1350 242
use SUNSAR_IVTRIX1_CV  XA3
timestamp 1708692311
transform 1 0 0 0 1 616
box -90 -66 1350 330
use SUNSAR_IVTRIX1_CV  XA4
timestamp 1708692311
transform 1 0 0 0 1 880
box -90 -66 1350 330
use SUNSAR_IVX1_CV  XA5
timestamp 1708692311
transform 1 0 0 0 1 1144
box -90 -66 1350 242
use SUNSAR_IVTRIX1_CV  XA6
timestamp 1708692311
transform 1 0 0 0 1 1320
box -90 -66 1350 330
use SUNSAR_NDTRIX1_CV  XA7
timestamp 1708692311
transform 1 0 0 0 1 1584
box -90 -66 1350 418
use SUNSAR_IVX1_CV  XA8
timestamp 1708692311
transform 1 0 0 0 1 1936
box -90 -66 1350 242
use SUNSAR_cut_M1M2_2x1  xcut0
timestamp 1708642800
transform 1 0 990 0 1 1039
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut1
timestamp 1708642800
transform 1 0 990 0 1 1479
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut2
timestamp 1708642800
transform 1 0 774 0 1 291
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut3
timestamp 1708642800
transform 1 0 162 0 1 775
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut4
timestamp 1708642800
transform 1 0 378 0 1 379
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut5
timestamp 1708642800
transform 1 0 162 0 1 1831
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut6
timestamp 1708642800
transform 1 0 990 0 1 1479
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut7
timestamp 1708642800
transform 1 0 378 0 1 1523
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut8
timestamp 1708642800
transform 1 0 378 0 1 1875
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut9
timestamp 1708642800
transform 1 0 162 0 1 1215
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut10
timestamp 1708642800
transform 1 0 378 0 1 1083
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut11
timestamp 1708642800
transform 1 0 774 0 1 1259
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut12
timestamp 1708642800
transform 1 0 990 0 1 951
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut13
timestamp 1708642800
transform 1 0 990 0 1 1391
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut14
timestamp 1708642800
transform 1 0 774 0 1 2051
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut15
timestamp 1708642800
transform 1 0 990 0 1 1743
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut16
timestamp 1708642800
transform 1 0 162 0 1 335
box 0 0 92 34
use SUNSAR_cut_M1M2_2x1  xcut17
timestamp 1708642800
transform 1 0 162 0 1 1655
box 0 0 92 34
<< labels >>
flabel locali s 162 687 270 721 0 FreeSans 200 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 200 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 378 2051 486 2085 0 FreeSans 200 0 0 0 Q
port 4 nsew signal bidirectional
flabel locali s 378 1875 486 1909 0 FreeSans 200 0 0 0 QN
port 5 nsew signal bidirectional
flabel locali s 162 1655 270 1689 0 FreeSans 200 0 0 0 RN
port 3 nsew signal bidirectional
flabel metal3 s 774 0 866 2112 0 FreeSans 200 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel metal3 s 378 0 470 2112 0 FreeSans 200 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 2112
<< end >>
