magic
tech sky130A
magscale 1 2
timestamp 1708902000
<< checkpaint >>
rect 0 0 1260 352
<< pdiff >>
rect 288 44 504 132
rect 288 132 504 220
rect 288 220 504 308
<< ntap >>
rect 1152 -44 1368 44
rect 1152 44 1368 132
rect 1152 132 1368 220
rect 1152 220 1368 308
rect 1152 308 1368 396
<< poly >>
rect 216 -18 936 18
rect 216 158 936 194
rect 216 334 936 370
rect 720 132 936 220
<< locali >>
rect 720 142 936 210
rect 1152 -44 1368 44
rect 288 54 504 122
rect 288 54 504 122
rect 1152 44 1368 132
rect 720 142 936 210
rect 1152 132 1368 220
rect 1152 132 1368 220
rect 288 230 504 298
rect 288 230 504 298
rect 1152 220 1368 308
rect 1152 308 1368 396
<< pcontact >>
rect 744 154 792 176
rect 744 176 792 198
rect 792 154 864 176
rect 792 176 864 198
rect 864 154 912 176
rect 864 176 912 198
<< ntapc >>
rect 1224 44 1296 132
rect 1224 220 1296 308
<< pdcontact >>
rect 312 66 360 88
rect 312 88 360 110
rect 360 66 432 88
rect 360 88 432 110
rect 432 66 480 88
rect 432 88 480 110
rect 312 242 360 264
rect 312 264 360 286
rect 360 242 432 264
rect 360 264 432 286
rect 432 242 480 264
rect 432 264 480 286
<< nwell >>
rect 0 -132 1440 484
<< labels >>
flabel locali s 720 142 936 210 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 54 504 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1152 132 1368 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 288 230 504 298 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 352
<< end >>
