magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 100 38
<< m3 >>
rect 0 0 100 38
<< v3 >>
rect 6 3 38 35
rect 62 3 94 35
<< m4 >>
rect 0 0 100 38
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 100 38
<< end >>
