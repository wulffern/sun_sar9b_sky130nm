magic
tech sky130A
magscale 1 2
timestamp 1708902000
<< checkpaint >>
rect 0 0 2520 528
<< poly >>
rect 324 158 2196 194
<< locali >>
rect 864 406 1032 474
rect 1032 54 1656 122
rect 1032 54 1100 474
rect 1656 54 1824 122
rect 1824 318 2088 386
rect 1824 54 1892 386
rect 830 230 898 298
rect 1622 230 1690 298
rect 2412 132 2628 220
rect -108 132 108 220
rect 1548 230 1764 298
rect 324 318 540 386
rect 1980 142 2196 210
rect 756 406 972 474
<< m3 >>
rect 1548 0 1732 528
rect 756 0 940 528
rect 1548 0 1732 528
rect 756 0 940 528
use SUNSAR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 176
box 0 176 1260 528
use SUNSAR_PCHDL MP0 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNSAR_PCHDL MP1 
transform 1 0 1260 0 1 176
box 1260 176 2520 528
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 406
box 1548 406 1732 474
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 756 0 1 54
box 756 54 940 122
<< labels >>
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 5 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 6 nsew signal bidirectional
flabel locali s 1548 230 1764 298 0 FreeSans 400 0 0 0 GNG
port 3 nsew signal bidirectional
flabel locali s 324 318 540 386 0 FreeSans 400 0 0 0 TIE_H
port 4 nsew signal bidirectional
flabel locali s 1980 142 2196 210 0 FreeSans 400 0 0 0 C
port 1 nsew signal bidirectional
flabel locali s 756 406 972 474 0 FreeSans 400 0 0 0 GN
port 2 nsew signal bidirectional
flabel m3 s 1548 0 1732 528 0 FreeSans 400 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel m3 s 756 0 940 528 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 528
<< end >>
