magic
tech sky130A
magscale 1 2
timestamp 1708642800
<< checkpaint >>
rect 0 0 68 184
<< m1 >>
rect 0 0 68 184
<< v1 >>
rect 6 12 62 68
rect 6 116 62 172
<< m2 >>
rect 0 0 68 184
<< v2 >>
rect 6 12 62 68
rect 6 116 62 172
<< m3 >>
rect 0 0 68 184
<< v3 >>
rect 6 12 62 68
rect 6 116 62 172
<< m4 >>
rect 0 0 68 184
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 68 184
<< end >>
