magic
tech sky130A
timestamp 1712959200
<< checkpaint >>
rect 0 0 34 96
<< metal3 >>
rect 0 90 34 92
rect 0 58 1 90
rect 33 58 34 90
rect 0 34 34 58
rect 0 2 1 34
rect 33 2 34 34
rect 0 0 34 2
<< via3 >>
rect 1 58 33 90
rect 1 2 33 34
<< metal4 >>
rect 0 90 34 96
rect 0 58 1 90
rect 33 58 34 90
rect 0 34 34 58
rect 0 2 1 34
rect 33 2 34 34
rect 0 0 34 2
<< properties >>
string FIXED_BBOX 0 0 34 96
<< end >>
