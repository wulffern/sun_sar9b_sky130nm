magic
tech sky130A
magscale 1 2
timestamp 1708902000
<< checkpaint >>
rect -2698 -1864 25806 51406
<< m3 >>
rect 8580 32744 23968 32812
rect 8580 33116 23968 33184
rect 23614 33456 23682 39884
rect 23890 33456 23958 44460
rect -690 33556 -622 43052
rect -690 33556 -622 43052
rect 3454 33742 3522 43052
rect 4350 33928 4418 43052
rect 8494 34114 8562 43052
rect 0 34300 68 43082
rect 2879 34486 2947 43082
rect 2879 34486 2947 43082
rect 5040 34672 5108 43082
rect 5040 34672 5108 43082
rect 7919 34858 7987 43082
rect 7919 34858 7987 43082
rect 10080 35044 10148 43082
rect 10080 35044 10148 43082
rect 12959 35230 13027 43082
rect 12959 35230 13027 43082
rect 15120 35416 15188 43082
rect 15120 35416 15188 43082
rect 17999 35602 18067 43082
rect 17999 35602 18067 43082
rect 143 35788 211 43962
rect 2736 35974 2804 43962
rect 5183 36160 5251 43962
rect 7776 36346 7844 43962
rect 300 36532 368 44842
rect 2580 36718 2648 44842
rect 5340 36904 5408 44842
rect 7620 37090 7688 44842
rect 10380 37276 10448 44842
rect 12660 37462 12728 44842
rect 15420 37648 15488 44842
rect 17700 37834 17768 44842
rect -290 38510 -106 49966
rect 3054 38510 3238 49966
rect 4750 38510 4934 49966
rect 8094 38510 8278 49966
rect 9790 38510 9974 49966
rect 13134 38510 13318 49966
rect 14830 38510 15014 49966
rect 18174 38510 18358 49966
rect 19870 38510 20054 49966
rect 23214 38510 23398 49966
rect 9174 -720 9358 4800
rect 13750 -720 13934 4800
rect 502 38510 686 50686
rect 2262 38510 2446 50686
rect 5542 38510 5726 50686
rect 7302 38510 7486 50686
rect 10582 38510 10766 50686
rect 12342 38510 12526 50686
rect 15622 38510 15806 50686
rect 17382 38510 17566 50686
rect 20662 38510 20846 50686
rect 22422 38510 22606 50686
rect 8382 -1440 8566 4800
rect 14542 -1440 14726 4800
rect 1078 42436 1262 51406
rect 1686 42436 1870 51406
rect 6118 42436 6302 51406
rect 6726 42436 6910 51406
rect 11158 42436 11342 51406
rect 11766 42436 11950 51406
rect 16198 42436 16382 51406
rect 16806 42436 16990 51406
rect 21238 42436 21422 51406
rect 9752 -1864 9820 2938
rect 13288 -1864 13356 2938
rect 10454 1110 10690 1178
rect 8614 4986 10454 5054
rect 12418 1110 12586 1178
rect 12586 4986 14494 5054
rect 10690 1110 10858 1178
rect 10858 2518 12418 2586
rect 10858 1110 10926 2586
rect 10582 230 10766 298
rect 12342 230 12526 298
rect 20160 43082 20228 43266
<< m2 >>
rect 14460 32254 14528 32812
rect 8580 32254 8648 33184
rect 23614 33116 23682 33456
rect 23890 32744 23958 33456
rect -690 33488 13976 33556
rect 3454 33674 13600 33742
rect 4350 33860 13224 33928
rect 8494 34046 12848 34114
rect 0 34232 9200 34300
rect 2879 34418 9576 34486
rect 5040 34604 9952 34672
rect 7919 34790 10328 34858
rect 10080 34976 10704 35044
rect 10824 35162 13027 35230
rect 11012 35348 15188 35416
rect 11200 35534 18067 35602
rect 143 35720 9388 35788
rect 2736 35906 9764 35974
rect 5183 36092 10140 36160
rect 7776 36278 10516 36346
rect 300 36464 13788 36532
rect 2580 36650 13412 36718
rect 5340 36836 13036 36904
rect 7620 37022 12660 37090
rect 10380 37208 12472 37276
rect 12216 37394 12728 37462
rect 12028 37580 15488 37648
rect 11840 37766 17768 37834
rect 502 48806 838 48874
rect 838 48204 3454 48272
rect 3386 48204 3454 48400
rect 838 48204 906 48874
rect 5542 48806 5878 48874
rect 5878 48204 8494 48272
rect 8426 48204 8494 48400
rect 5878 48204 5946 48874
rect 10582 48806 10918 48874
rect 10918 48204 13534 48272
rect 13466 48204 13534 48400
rect 10918 48204 10986 48874
rect 15622 48806 15958 48874
rect 15958 48204 18574 48272
rect 18506 48204 18574 48400
rect 15958 48204 16026 48874
rect -722 45740 19654 45808
rect -790 45740 -722 45936
rect 3386 45740 3454 45936
rect 4250 45740 4318 45936
rect 8426 45740 8494 45936
rect 9290 45740 9358 45936
rect 13466 45740 13534 45936
rect 14330 45740 14398 45936
rect 18506 45740 18574 45936
rect 19370 45740 19438 45936
rect 534 39268 838 39336
rect 838 38876 3454 38944
rect 3386 38876 3454 39072
rect 838 38876 906 39336
rect 5574 39268 5878 39336
rect 5878 38876 8494 38944
rect 8426 38876 8494 39072
rect 5878 38876 5946 39336
rect 10614 39268 10918 39336
rect 10918 38876 13534 38944
rect 13466 38876 13534 39072
rect 10918 38876 10986 39336
rect 15654 39268 15958 39336
rect 15958 38876 18574 38944
rect 18506 38876 18574 39072
rect 15958 38876 16026 39336
rect 20694 39268 20998 39336
rect 20998 39268 21066 39336
rect 2230 39268 2534 39336
rect 2534 39268 2602 39396
rect 2534 39396 4350 39464
rect 4282 39004 4350 39464
rect 7270 39268 7574 39336
rect 7574 39268 7642 39396
rect 7574 39396 9390 39464
rect 9322 39004 9390 39464
rect 12310 39268 12614 39336
rect 12614 39268 12682 39396
rect 12614 39396 14430 39464
rect 14362 39004 14430 39464
rect 17350 39268 17654 39336
rect 17654 39268 17722 39396
rect 17654 39396 19470 39464
rect 19402 39004 19470 39464
rect -690 41040 19654 41108
rect -758 40764 -690 41108
rect 3386 40764 3454 41108
rect 4282 40764 4350 41108
rect 8426 40764 8494 41108
rect 9322 40764 9390 41108
rect 13466 40764 13534 41108
rect 14362 40764 14430 41108
rect 18506 40764 18574 41108
rect 19402 40764 19470 41108
rect -722 41192 19654 41260
rect -790 41192 -722 41536
rect 3386 41192 3454 41536
rect 4250 41192 4318 41536
rect 8426 41192 8494 41536
rect 9290 41192 9358 41536
rect 13466 41192 13534 41536
rect 14330 41192 14398 41536
rect 18506 41192 18574 41536
rect 19370 41192 19438 41536
rect -506 41820 934 41888
rect 934 41820 2014 41888
rect 934 41820 6190 41888
rect 934 41820 7054 41888
rect 934 41820 11230 41888
rect 934 41820 12094 41888
rect 934 41820 16270 41888
rect 934 41820 17134 41888
rect 934 41820 21310 41888
rect 22922 41942 23290 42010
rect 19594 40832 22922 40900
rect 22922 40832 22990 42010
rect 19562 40764 19654 40832
rect 22262 42822 22498 42890
rect 19594 41536 22262 41604
rect 22262 41536 22330 42890
rect 19546 41468 19654 41536
rect 22066 47276 22234 47344
rect 19546 46220 22234 46288
rect 22234 46220 22302 47344
rect 21830 47804 22066 47872
rect 20770 48806 21830 48874
rect 21830 47804 21898 48874
rect 10690 2518 10858 2586
rect 10858 1110 12418 1178
rect 10858 1110 10926 2586
rect -722 41820 1150 41888
<< m1 >>
rect 13908 32186 13976 33488
rect 13532 32186 13600 33674
rect 13156 32186 13224 33860
rect 12780 32186 12848 34046
rect 9132 32186 9200 34232
rect 9508 32186 9576 34418
rect 9884 32186 9952 34604
rect 10260 32186 10328 34790
rect 10636 32186 10704 34976
rect 10824 32186 10892 35162
rect 11012 32186 11080 35348
rect 11200 32186 11268 35534
rect 9320 32186 9388 35720
rect 9696 32186 9764 35906
rect 10072 32186 10140 36092
rect 10448 32186 10516 36278
rect 13720 32186 13788 36464
rect 13344 32186 13412 36650
rect 12968 32186 13036 36836
rect 12592 32186 12660 37022
rect 12404 32186 12472 37208
rect 12216 32186 12284 37394
rect 12028 32186 12096 37580
rect 11840 32186 11908 37766
rect 9648 -1652 9716 562
rect 13392 -1652 13460 562
rect -2630 48332 -722 48400
rect 2230 48772 2566 48840
rect 2566 48204 4318 48272
rect 4250 48204 4318 48400
rect 2566 48204 2634 48840
rect 7270 48772 7606 48840
rect 7606 48204 9358 48272
rect 9290 48204 9358 48400
rect 7606 48204 7674 48840
rect 12310 48772 12646 48840
rect 12646 48204 14398 48272
rect 14330 48204 14398 48400
rect 12646 48204 12714 48840
rect 17350 48772 17686 48840
rect 17686 48204 19438 48272
rect 19370 48204 19438 48400
rect 17686 48204 17754 48840
rect 21830 47452 22066 47520
rect 19978 47012 21830 47080
rect 21830 47012 21898 47520
rect -1766 4986 68 5054
rect -1766 8386 68 8454
rect -1766 11786 68 11854
rect -1766 15186 68 15254
rect -1766 18586 68 18654
rect -1766 21986 68 22054
rect -1766 25386 68 25454
rect -1766 28786 68 28854
rect 23040 4986 24874 5054
rect 23040 8386 24874 8454
rect 23040 11786 24874 11854
rect 23040 15186 24874 15254
rect 23040 18586 24874 18654
rect 23040 21986 24874 22054
rect 23040 25386 24874 25454
rect 23040 28786 24874 28854
<< locali >>
rect 24690 -720 24874 49966
rect -1766 -720 24874 -536
rect -1766 49782 24874 49966
rect -1766 -720 -1582 49966
rect 24690 -720 24874 49966
rect 25410 -1440 25594 50686
rect -2486 -1440 25594 -1256
rect -2486 50502 25594 50686
rect -2486 -1440 -2302 50686
rect 25410 -1440 25594 50686
rect -2486 51222 25594 51406
rect -2486 51222 25594 51406
rect 25738 -1652 25806 51406
rect -2486 -1652 25806 -1584
rect 25738 -1652 25806 51406
rect -2698 -1864 25806 -1796
rect -2698 -1864 -2630 51406
rect 19870 47012 20086 47080
rect -722 45868 -506 45936
rect 934 41820 1150 41888
rect 10582 2518 10798 2586
rect 10582 1110 10798 1178
<< m4 >>
rect 10454 1110 10522 5054
rect 12586 1110 12654 5054
use SUNSAR_SARBSSW_CV XB1 
transform -1 0 11554 0 1 0
box 11554 0 23002 4800
use SUNSAR_SARBSSW_CV XB2 
transform 1 0 11554 0 1 0
box 11554 0 23002 4800
use SUNSAR_CDAC8_CV XDAC1 
transform -1 0 11404 0 1 4986
box 11404 4986 22672 32254
use SUNSAR_CDAC8_CV XDAC2 
transform 1 0 11704 0 1 4986
box 11704 4986 22972 32254
use SUNSAR_SARDIGEX4_CV XA0 
transform 1 0 -1046 0 1 38510
box -1046 38510 1474 49246
use SUNSAR_SARDIGEX4_CV XA1 
transform -1 0 3994 0 1 38510
box 3994 38510 6514 49246
use SUNSAR_SARDIGEX4_CV XA2 
transform 1 0 3994 0 1 38510
box 3994 38510 6514 49246
use SUNSAR_SARDIGEX4_CV XA3 
transform -1 0 9034 0 1 38510
box 9034 38510 11554 49246
use SUNSAR_SARDIGEX4_CV XA4 
transform 1 0 9034 0 1 38510
box 9034 38510 11554 49246
use SUNSAR_SARDIGEX4_CV XA5 
transform -1 0 14074 0 1 38510
box 14074 38510 16594 49246
use SUNSAR_SARDIGEX4_CV XA6 
transform 1 0 14074 0 1 38510
box 14074 38510 16594 49246
use SUNSAR_SARDIGEX4_CV XA7 
transform -1 0 19114 0 1 38510
box 19114 38510 21634 49246
use SUNSAR_SARDIGEX4_CV XA8 
transform 1 0 19114 0 1 38510
box 19114 38510 21634 49246
use SUNSAR_SARCMPX1_CV XA20 
transform -1 0 24154 0 1 38510
box 24154 38510 26674 48366
use SUNSAR_cut_M3M4_1x2 xcut0 
transform 1 0 14460 0 1 32254
box 14460 32254 14528 32438
use SUNSAR_cut_M3M4_2x1 xcut1 
transform 1 0 14460 0 1 32744
box 14460 32744 14644 32812
use SUNSAR_cut_M3M4_1x2 xcut2 
transform 1 0 8580 0 1 32254
box 8580 32254 8648 32438
use SUNSAR_cut_M3M4_2x1 xcut3 
transform 1 0 8580 0 1 33116
box 8580 33116 8764 33184
use SUNSAR_cut_M2M4_2x1 xcut4 
transform 1 0 23614 0 1 39884
box 23614 39884 23798 39952
use SUNSAR_cut_M3M4_2x1 xcut5 
transform 1 0 23614 0 1 33116
box 23614 33116 23798 33184
use SUNSAR_cut_M3M4_1x2 xcut6 
transform 1 0 23614 0 1 33456
box 23614 33456 23682 33640
use SUNSAR_cut_M3M4_2x1 xcut7 
transform 1 0 23774 0 1 44460
box 23774 44460 23958 44528
use SUNSAR_cut_M2M3_2x1 xcut8 
transform 1 0 23614 0 1 44460
box 23614 44460 23798 44528
use SUNSAR_cut_M3M4_2x1 xcut9 
transform 1 0 23890 0 1 32744
box 23890 32744 24074 32812
use SUNSAR_cut_M3M4_1x2 xcut10 
transform 1 0 23890 0 1 33456
box 23890 33456 23958 33640
use SUNSAR_cut_M3M4_1x2 xcut11 
transform 1 0 -690 0 1 33430
box -690 33430 -622 33614
use SUNSAR_cut_M2M3_1x2 xcut12 
transform 1 0 13908 0 1 33430
box 13908 33430 13976 33614
use SUNSAR_cut_M3M4_1x2 xcut13 
transform 1 0 3454 0 1 33616
box 3454 33616 3522 33800
use SUNSAR_cut_M2M3_1x2 xcut14 
transform 1 0 13532 0 1 33616
box 13532 33616 13600 33800
use SUNSAR_cut_M3M4_1x2 xcut15 
transform 1 0 4350 0 1 33802
box 4350 33802 4418 33986
use SUNSAR_cut_M2M3_1x2 xcut16 
transform 1 0 13156 0 1 33802
box 13156 33802 13224 33986
use SUNSAR_cut_M3M4_1x2 xcut17 
transform 1 0 8494 0 1 33988
box 8494 33988 8562 34172
use SUNSAR_cut_M2M3_1x2 xcut18 
transform 1 0 12780 0 1 33988
box 12780 33988 12848 34172
use SUNSAR_cut_M3M4_1x2 xcut19 
transform 1 0 0 0 1 34174
box 0 34174 68 34358
use SUNSAR_cut_M2M3_1x2 xcut20 
transform 1 0 9132 0 1 34174
box 9132 34174 9200 34358
use SUNSAR_cut_M3M4_1x2 xcut21 
transform 1 0 2879 0 1 34360
box 2879 34360 2947 34544
use SUNSAR_cut_M2M3_1x2 xcut22 
transform 1 0 9508 0 1 34360
box 9508 34360 9576 34544
use SUNSAR_cut_M3M4_1x2 xcut23 
transform 1 0 5040 0 1 34546
box 5040 34546 5108 34730
use SUNSAR_cut_M2M3_1x2 xcut24 
transform 1 0 9884 0 1 34546
box 9884 34546 9952 34730
use SUNSAR_cut_M3M4_1x2 xcut25 
transform 1 0 7919 0 1 34732
box 7919 34732 7987 34916
use SUNSAR_cut_M2M3_1x2 xcut26 
transform 1 0 10260 0 1 34732
box 10260 34732 10328 34916
use SUNSAR_cut_M3M4_1x2 xcut27 
transform 1 0 10080 0 1 34918
box 10080 34918 10148 35102
use SUNSAR_cut_M2M3_1x2 xcut28 
transform 1 0 10636 0 1 34918
box 10636 34918 10704 35102
use SUNSAR_cut_M3M4_1x2 xcut29 
transform 1 0 12959 0 1 35104
box 12959 35104 13027 35288
use SUNSAR_cut_M2M3_1x2 xcut30 
transform 1 0 10824 0 1 35104
box 10824 35104 10892 35288
use SUNSAR_cut_M3M4_1x2 xcut31 
transform 1 0 15120 0 1 35290
box 15120 35290 15188 35474
use SUNSAR_cut_M2M3_1x2 xcut32 
transform 1 0 11012 0 1 35290
box 11012 35290 11080 35474
use SUNSAR_cut_M3M4_1x2 xcut33 
transform 1 0 17999 0 1 35476
box 17999 35476 18067 35660
use SUNSAR_cut_M2M3_1x2 xcut34 
transform 1 0 11200 0 1 35476
box 11200 35476 11268 35660
use SUNSAR_cut_M3M4_1x2 xcut35 
transform 1 0 143 0 1 35662
box 143 35662 211 35846
use SUNSAR_cut_M2M3_1x2 xcut36 
transform 1 0 9320 0 1 35662
box 9320 35662 9388 35846
use SUNSAR_cut_M3M4_1x2 xcut37 
transform 1 0 2736 0 1 35848
box 2736 35848 2804 36032
use SUNSAR_cut_M2M3_1x2 xcut38 
transform 1 0 9696 0 1 35848
box 9696 35848 9764 36032
use SUNSAR_cut_M3M4_1x2 xcut39 
transform 1 0 5183 0 1 36034
box 5183 36034 5251 36218
use SUNSAR_cut_M2M3_1x2 xcut40 
transform 1 0 10072 0 1 36034
box 10072 36034 10140 36218
use SUNSAR_cut_M3M4_1x2 xcut41 
transform 1 0 7776 0 1 36220
box 7776 36220 7844 36404
use SUNSAR_cut_M2M3_1x2 xcut42 
transform 1 0 10448 0 1 36220
box 10448 36220 10516 36404
use SUNSAR_cut_M3M4_1x2 xcut43 
transform 1 0 300 0 1 36406
box 300 36406 368 36590
use SUNSAR_cut_M2M3_1x2 xcut44 
transform 1 0 13720 0 1 36406
box 13720 36406 13788 36590
use SUNSAR_cut_M3M4_1x2 xcut45 
transform 1 0 2580 0 1 36592
box 2580 36592 2648 36776
use SUNSAR_cut_M2M3_1x2 xcut46 
transform 1 0 13344 0 1 36592
box 13344 36592 13412 36776
use SUNSAR_cut_M3M4_1x2 xcut47 
transform 1 0 5340 0 1 36778
box 5340 36778 5408 36962
use SUNSAR_cut_M2M3_1x2 xcut48 
transform 1 0 12968 0 1 36778
box 12968 36778 13036 36962
use SUNSAR_cut_M3M4_1x2 xcut49 
transform 1 0 7620 0 1 36964
box 7620 36964 7688 37148
use SUNSAR_cut_M2M3_1x2 xcut50 
transform 1 0 12592 0 1 36964
box 12592 36964 12660 37148
use SUNSAR_cut_M3M4_1x2 xcut51 
transform 1 0 10380 0 1 37150
box 10380 37150 10448 37334
use SUNSAR_cut_M2M3_1x2 xcut52 
transform 1 0 12404 0 1 37150
box 12404 37150 12472 37334
use SUNSAR_cut_M3M4_1x2 xcut53 
transform 1 0 12660 0 1 37336
box 12660 37336 12728 37520
use SUNSAR_cut_M2M3_1x2 xcut54 
transform 1 0 12216 0 1 37336
box 12216 37336 12284 37520
use SUNSAR_cut_M3M4_1x2 xcut55 
transform 1 0 15420 0 1 37522
box 15420 37522 15488 37706
use SUNSAR_cut_M2M3_1x2 xcut56 
transform 1 0 12028 0 1 37522
box 12028 37522 12096 37706
use SUNSAR_cut_M3M4_1x2 xcut57 
transform 1 0 17700 0 1 37708
box 17700 37708 17768 37892
use SUNSAR_cut_M2M3_1x2 xcut58 
transform 1 0 11840 0 1 37708
box 11840 37708 11908 37892
use SUNSAR_cut_M1M4_2x2 xcut59 
transform 1 0 -290 0 1 49782
box -290 49782 -106 49966
use SUNSAR_cut_M1M4_2x2 xcut60 
transform 1 0 3054 0 1 49782
box 3054 49782 3238 49966
use SUNSAR_cut_M1M4_2x2 xcut61 
transform 1 0 4750 0 1 49782
box 4750 49782 4934 49966
use SUNSAR_cut_M1M4_2x2 xcut62 
transform 1 0 8094 0 1 49782
box 8094 49782 8278 49966
use SUNSAR_cut_M1M4_2x2 xcut63 
transform 1 0 9790 0 1 49782
box 9790 49782 9974 49966
use SUNSAR_cut_M1M4_2x2 xcut64 
transform 1 0 13134 0 1 49782
box 13134 49782 13318 49966
use SUNSAR_cut_M1M4_2x2 xcut65 
transform 1 0 14830 0 1 49782
box 14830 49782 15014 49966
use SUNSAR_cut_M1M4_2x2 xcut66 
transform 1 0 18174 0 1 49782
box 18174 49782 18358 49966
use SUNSAR_cut_M1M4_2x2 xcut67 
transform 1 0 19870 0 1 49782
box 19870 49782 20054 49966
use SUNSAR_cut_M1M4_2x2 xcut68 
transform 1 0 23214 0 1 49782
box 23214 49782 23398 49966
use SUNSAR_cut_M1M4_2x2 xcut69 
transform 1 0 9174 0 1 -720
box 9174 -720 9358 -536
use SUNSAR_cut_M1M4_2x2 xcut70 
transform 1 0 13750 0 1 -720
box 13750 -720 13934 -536
use SUNSAR_cut_M1M4_2x2 xcut71 
transform 1 0 502 0 1 50502
box 502 50502 686 50686
use SUNSAR_cut_M1M4_2x2 xcut72 
transform 1 0 2262 0 1 50502
box 2262 50502 2446 50686
use SUNSAR_cut_M1M4_2x2 xcut73 
transform 1 0 5542 0 1 50502
box 5542 50502 5726 50686
use SUNSAR_cut_M1M4_2x2 xcut74 
transform 1 0 7302 0 1 50502
box 7302 50502 7486 50686
use SUNSAR_cut_M1M4_2x2 xcut75 
transform 1 0 10582 0 1 50502
box 10582 50502 10766 50686
use SUNSAR_cut_M1M4_2x2 xcut76 
transform 1 0 12342 0 1 50502
box 12342 50502 12526 50686
use SUNSAR_cut_M1M4_2x2 xcut77 
transform 1 0 15622 0 1 50502
box 15622 50502 15806 50686
use SUNSAR_cut_M1M4_2x2 xcut78 
transform 1 0 17382 0 1 50502
box 17382 50502 17566 50686
use SUNSAR_cut_M1M4_2x2 xcut79 
transform 1 0 20662 0 1 50502
box 20662 50502 20846 50686
use SUNSAR_cut_M1M4_2x2 xcut80 
transform 1 0 22422 0 1 50502
box 22422 50502 22606 50686
use SUNSAR_cut_M1M4_2x2 xcut81 
transform 1 0 8382 0 1 -1440
box 8382 -1440 8566 -1256
use SUNSAR_cut_M1M4_2x2 xcut82 
transform 1 0 14542 0 1 -1440
box 14542 -1440 14726 -1256
use SUNSAR_cut_M1M4_2x2 xcut83 
transform 1 0 1078 0 1 51222
box 1078 51222 1262 51406
use SUNSAR_cut_M1M4_2x2 xcut84 
transform 1 0 1686 0 1 51222
box 1686 51222 1870 51406
use SUNSAR_cut_M1M4_2x2 xcut85 
transform 1 0 6118 0 1 51222
box 6118 51222 6302 51406
use SUNSAR_cut_M1M4_2x2 xcut86 
transform 1 0 6726 0 1 51222
box 6726 51222 6910 51406
use SUNSAR_cut_M1M4_2x2 xcut87 
transform 1 0 11158 0 1 51222
box 11158 51222 11342 51406
use SUNSAR_cut_M1M4_2x2 xcut88 
transform 1 0 11766 0 1 51222
box 11766 51222 11950 51406
use SUNSAR_cut_M1M4_2x2 xcut89 
transform 1 0 16198 0 1 51222
box 16198 51222 16382 51406
use SUNSAR_cut_M1M4_2x2 xcut90 
transform 1 0 16806 0 1 51222
box 16806 51222 16990 51406
use SUNSAR_cut_M1M4_2x2 xcut91 
transform 1 0 21238 0 1 51222
box 21238 51222 21422 51406
use SUNSAR_cut_M1M2_2x1 xcut92 
transform 1 0 9590 0 1 494
box 9590 494 9774 562
use SUNSAR_cut_M1M2_2x1 xcut93 
transform 1 0 9590 0 1 -1652
box 9590 -1652 9774 -1584
use SUNSAR_cut_M1M2_2x1 xcut94 
transform 1 0 13334 0 1 494
box 13334 494 13518 562
use SUNSAR_cut_M1M2_2x1 xcut95 
transform 1 0 13334 0 1 -1652
box 13334 -1652 13518 -1584
use SUNSAR_cut_M1M2_2x1 xcut96 
transform 1 0 -722 0 1 48332
box -722 48332 -538 48400
use SUNSAR_cut_M1M2_1x2 xcut97 
transform 1 0 -2698 0 1 48274
box -2698 48274 -2630 48458
use SUNSAR_cut_M1M4_2x1 xcut98 
transform 1 0 9694 0 1 -1864
box 9694 -1864 9878 -1796
use SUNSAR_cut_M1M4_2x1 xcut99 
transform 1 0 13230 0 1 -1864
box 13230 -1864 13414 -1796
use SUNSAR_cut_M1M3_2x1 xcut100 
transform 1 0 502 0 1 48806
box 502 48806 686 48874
use SUNSAR_cut_M1M3_2x1 xcut101 
transform 1 0 3454 0 1 48332
box 3454 48332 3638 48400
use SUNSAR_cut_M1M3_2x1 xcut102 
transform 1 0 5542 0 1 48806
box 5542 48806 5726 48874
use SUNSAR_cut_M1M3_2x1 xcut103 
transform 1 0 8494 0 1 48332
box 8494 48332 8678 48400
use SUNSAR_cut_M1M3_2x1 xcut104 
transform 1 0 10582 0 1 48806
box 10582 48806 10766 48874
use SUNSAR_cut_M1M3_2x1 xcut105 
transform 1 0 13534 0 1 48332
box 13534 48332 13718 48400
use SUNSAR_cut_M1M3_2x1 xcut106 
transform 1 0 15622 0 1 48806
box 15622 48806 15806 48874
use SUNSAR_cut_M1M3_2x1 xcut107 
transform 1 0 18574 0 1 48332
box 18574 48332 18758 48400
use SUNSAR_cut_M1M3_2x1 xcut108 
transform 1 0 -722 0 1 45868
box -722 45868 -538 45936
use SUNSAR_cut_M1M3_2x1 xcut109 
transform 1 0 3454 0 1 45868
box 3454 45868 3638 45936
use SUNSAR_cut_M1M3_2x1 xcut110 
transform 1 0 4318 0 1 45868
box 4318 45868 4502 45936
use SUNSAR_cut_M1M3_2x1 xcut111 
transform 1 0 8494 0 1 45868
box 8494 45868 8678 45936
use SUNSAR_cut_M1M3_2x1 xcut112 
transform 1 0 9358 0 1 45868
box 9358 45868 9542 45936
use SUNSAR_cut_M1M3_2x1 xcut113 
transform 1 0 13534 0 1 45868
box 13534 45868 13718 45936
use SUNSAR_cut_M1M3_2x1 xcut114 
transform 1 0 14398 0 1 45868
box 14398 45868 14582 45936
use SUNSAR_cut_M1M3_2x1 xcut115 
transform 1 0 18574 0 1 45868
box 18574 45868 18758 45936
use SUNSAR_cut_M1M3_2x1 xcut116 
transform 1 0 19438 0 1 45868
box 19438 45868 19622 45936
use SUNSAR_cut_M1M2_2x1 xcut117 
transform 1 0 2230 0 1 48772
box 2230 48772 2414 48840
use SUNSAR_cut_M1M2_2x1 xcut118 
transform 1 0 4318 0 1 48332
box 4318 48332 4502 48400
use SUNSAR_cut_M1M2_2x1 xcut119 
transform 1 0 7270 0 1 48772
box 7270 48772 7454 48840
use SUNSAR_cut_M1M2_2x1 xcut120 
transform 1 0 9358 0 1 48332
box 9358 48332 9542 48400
use SUNSAR_cut_M1M2_2x1 xcut121 
transform 1 0 12310 0 1 48772
box 12310 48772 12494 48840
use SUNSAR_cut_M1M2_2x1 xcut122 
transform 1 0 14398 0 1 48332
box 14398 48332 14582 48400
use SUNSAR_cut_M1M2_2x1 xcut123 
transform 1 0 17350 0 1 48772
box 17350 48772 17534 48840
use SUNSAR_cut_M1M2_2x1 xcut124 
transform 1 0 19438 0 1 48332
box 19438 48332 19622 48400
use SUNSAR_cut_M1M3_2x1 xcut125 
transform 1 0 -722 0 1 41468
box -722 41468 -538 41536
use SUNSAR_cut_M1M3_2x1 xcut126 
transform 1 0 3454 0 1 41468
box 3454 41468 3638 41536
use SUNSAR_cut_M1M3_2x1 xcut127 
transform 1 0 4318 0 1 41468
box 4318 41468 4502 41536
use SUNSAR_cut_M1M3_2x1 xcut128 
transform 1 0 8494 0 1 41468
box 8494 41468 8678 41536
use SUNSAR_cut_M1M3_2x1 xcut129 
transform 1 0 9358 0 1 41468
box 9358 41468 9542 41536
use SUNSAR_cut_M1M3_2x1 xcut130 
transform 1 0 13534 0 1 41468
box 13534 41468 13718 41536
use SUNSAR_cut_M1M3_2x1 xcut131 
transform 1 0 14398 0 1 41468
box 14398 41468 14582 41536
use SUNSAR_cut_M1M3_2x1 xcut132 
transform 1 0 18574 0 1 41468
box 18574 41468 18758 41536
use SUNSAR_cut_M1M3_2x1 xcut133 
transform 1 0 19438 0 1 41468
box 19438 41468 19622 41536
use SUNSAR_cut_M1M3_2x1 xcut134 
transform 1 0 934 0 1 41820
box 934 41820 1118 41888
use SUNSAR_cut_M1M3_2x1 xcut135 
transform 1 0 1798 0 1 41820
box 1798 41820 1982 41888
use SUNSAR_cut_M1M3_2x1 xcut136 
transform 1 0 5974 0 1 41820
box 5974 41820 6158 41888
use SUNSAR_cut_M1M3_2x1 xcut137 
transform 1 0 6838 0 1 41820
box 6838 41820 7022 41888
use SUNSAR_cut_M1M3_2x1 xcut138 
transform 1 0 11014 0 1 41820
box 11014 41820 11198 41888
use SUNSAR_cut_M1M3_2x1 xcut139 
transform 1 0 11878 0 1 41820
box 11878 41820 12062 41888
use SUNSAR_cut_M1M3_2x1 xcut140 
transform 1 0 16054 0 1 41820
box 16054 41820 16238 41888
use SUNSAR_cut_M1M3_2x1 xcut141 
transform 1 0 16918 0 1 41820
box 16918 41820 17102 41888
use SUNSAR_cut_M1M3_2x1 xcut142 
transform 1 0 21094 0 1 41820
box 21094 41820 21278 41888
use SUNSAR_cut_M1M3_2x1 xcut143 
transform 1 0 23214 0 1 41942
box 23214 41942 23398 42010
use SUNSAR_cut_M1M3_2x1 xcut144 
transform 1 0 22422 0 1 42822
box 22422 42822 22606 42890
use SUNSAR_cut_M1M3_2x1 xcut145 
transform 1 0 21958 0 1 47276
box 21958 47276 22142 47344
use SUNSAR_cut_M1M3_2x1 xcut146 
transform 1 0 19438 0 1 46220
box 19438 46220 19622 46288
use SUNSAR_cut_M1M3_2x1 xcut147 
transform 1 0 21990 0 1 47804
box 21990 47804 22174 47872
use SUNSAR_cut_M1M3_2x1 xcut148 
transform 1 0 20694 0 1 48806
box 20694 48806 20878 48874
use SUNSAR_cut_M1M2_2x1 xcut149 
transform 1 0 21990 0 1 47452
box 21990 47452 22174 47520
use SUNSAR_cut_M1M2_2x1 xcut150 
transform 1 0 19902 0 1 47012
box 19902 47012 20086 47080
use SUNSAR_cut_M4M5_1x2 xcut151 
transform 1 0 10454 0 1 1110
box 10454 1110 10522 1294
use SUNSAR_cut_M4M5_1x2 xcut152 
transform 1 0 10454 0 1 4870
box 10454 4870 10522 5054
use SUNSAR_cut_M1M4_2x1 xcut153 
transform 1 0 12310 0 1 1110
box 12310 1110 12494 1178
use SUNSAR_cut_M4M5_1x2 xcut154 
transform 1 0 12586 0 1 1110
box 12586 1110 12654 1294
use SUNSAR_cut_M4M5_1x2 xcut155 
transform 1 0 12586 0 1 4870
box 12586 4870 12654 5054
use SUNSAR_cut_M1M3_2x1 xcut156 
transform 1 0 10582 0 1 2518
box 10582 2518 10766 2586
use SUNSAR_cut_M1M3_2x1 xcut157 
transform 1 0 12310 0 1 1110
box 12310 1110 12494 1178
use SUNSAR_cut_M1M4_2x1 xcut158 
transform 1 0 10582 0 1 1110
box 10582 1110 10766 1178
use SUNSAR_cut_M1M4_2x1 xcut159 
transform 1 0 12310 0 1 2518
box 12310 2518 12494 2586
use SUNSAR_cut_M1M3_2x1 xcut160 
transform 1 0 -722 0 1 41820
box -722 41820 -538 41888
use SUNSAR_cut_M1M2_2x2 xcut161 
transform 1 0 -1766 0 1 5054
box -1766 5054 -1582 5238
use SUNSAR_cut_M1M2_2x2 xcut162 
transform 1 0 -1766 0 1 8454
box -1766 8454 -1582 8638
use SUNSAR_cut_M1M2_2x2 xcut163 
transform 1 0 -1766 0 1 11854
box -1766 11854 -1582 12038
use SUNSAR_cut_M1M2_2x2 xcut164 
transform 1 0 -1766 0 1 15254
box -1766 15254 -1582 15438
use SUNSAR_cut_M1M2_2x2 xcut165 
transform 1 0 -1766 0 1 18654
box -1766 18654 -1582 18838
use SUNSAR_cut_M1M2_2x2 xcut166 
transform 1 0 -1766 0 1 22054
box -1766 22054 -1582 22238
use SUNSAR_cut_M1M2_2x2 xcut167 
transform 1 0 -1766 0 1 25454
box -1766 25454 -1582 25638
use SUNSAR_cut_M1M2_2x2 xcut168 
transform 1 0 -1766 0 1 28854
box -1766 28854 -1582 29038
use SUNSAR_cut_M1M2_1x2 xcut169 
transform 1 0 24806 0 1 4986
box 24806 4986 24874 5170
use SUNSAR_cut_M1M2_1x2 xcut170 
transform 1 0 24806 0 1 8386
box 24806 8386 24874 8570
use SUNSAR_cut_M1M2_1x2 xcut171 
transform 1 0 24806 0 1 11786
box 24806 11786 24874 11970
use SUNSAR_cut_M1M2_1x2 xcut172 
transform 1 0 24806 0 1 15186
box 24806 15186 24874 15370
use SUNSAR_cut_M1M2_1x2 xcut173 
transform 1 0 24806 0 1 18586
box 24806 18586 24874 18770
use SUNSAR_cut_M1M2_1x2 xcut174 
transform 1 0 24806 0 1 21986
box 24806 21986 24874 22170
use SUNSAR_cut_M1M2_1x2 xcut175 
transform 1 0 24806 0 1 25386
box 24806 25386 24874 25570
use SUNSAR_cut_M1M2_1x2 xcut176 
transform 1 0 24806 0 1 28786
box 24806 28786 24874 28970
<< labels >>
flabel m3 s -690 33556 -622 43052 0 FreeSans 400 0 0 0 D<8>
port 6 nsew signal bidirectional
flabel m3 s 2879 34486 2947 43082 0 FreeSans 400 0 0 0 D<7>
port 7 nsew signal bidirectional
flabel m3 s 5040 34672 5108 43082 0 FreeSans 400 0 0 0 D<6>
port 8 nsew signal bidirectional
flabel m3 s 7919 34858 7987 43082 0 FreeSans 400 0 0 0 D<5>
port 9 nsew signal bidirectional
flabel m3 s 10080 35044 10148 43082 0 FreeSans 400 0 0 0 D<4>
port 10 nsew signal bidirectional
flabel m3 s 12959 35230 13027 43082 0 FreeSans 400 0 0 0 D<3>
port 11 nsew signal bidirectional
flabel m3 s 15120 35416 15188 43082 0 FreeSans 400 0 0 0 D<2>
port 12 nsew signal bidirectional
flabel m3 s 17999 35602 18067 43082 0 FreeSans 400 0 0 0 D<1>
port 13 nsew signal bidirectional
flabel locali s 24690 -720 24874 49966 0 FreeSans 400 0 0 0 AVSS
port 20 nsew signal bidirectional
flabel locali s 25410 -1440 25594 50686 0 FreeSans 400 0 0 0 AVDD
port 19 nsew signal bidirectional
flabel locali s -2486 51222 25594 51406 0 FreeSans 400 0 0 0 VREF
port 18 nsew signal bidirectional
flabel locali s 25738 -1652 25806 51406 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew signal bidirectional
flabel locali s 19870 47012 20086 47080 0 FreeSans 400 0 0 0 DONE
port 5 nsew signal bidirectional
flabel m3 s 10582 230 10766 298 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew signal bidirectional
flabel m3 s 12342 230 12526 298 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew signal bidirectional
flabel locali s -722 45868 -506 45936 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew signal bidirectional
flabel locali s 934 41820 1150 41888 0 FreeSans 400 0 0 0 EN
port 15 nsew signal bidirectional
flabel locali s 10582 2518 10798 2586 0 FreeSans 400 0 0 0 SARN
port 3 nsew signal bidirectional
flabel locali s 10582 1110 10798 1178 0 FreeSans 400 0 0 0 SARP
port 4 nsew signal bidirectional
flabel m3 s 20160 43082 20228 43266 0 FreeSans 400 0 0 0 D<0>
port 14 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -2698 -1864 25806 51406
<< end >>
