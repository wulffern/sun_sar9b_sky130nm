magic
tech sky130B
timestamp 1681336800
<< locali >>
rect 0 0 30 38
rect 60 0 90 38
<< rlocali >>
rect 30 0 60 38
<< labels >>
flabel locali s 0 0 30 38 0 FreeSans 200 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 30 0 90 38 0 FreeSans 200 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 60 0
<< end >>
