magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 1260 176
<< locali >>
rect -54 71 270 105
rect 216 71 300 105
rect 300 27 432 61
rect 300 27 334 105
rect 216 71 300 105
rect 300 115 432 149
rect 300 71 334 149
rect 828 27 912 61
rect 912 71 1044 105
rect 912 27 946 105
rect 828 115 912 149
rect 912 71 1044 105
rect 912 71 946 149
rect 990 71 1314 105
<< m3 >>
rect 774 0 874 176
rect 378 0 478 176
rect 774 0 874 176
rect 378 0 478 176
use SUNSAR_NCHDL MN1 
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNSAR_PCHDL MP1 
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNSAR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 115
box 774 115 874 153
use SUNSAR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 27
box 774 27 874 65
use SUNSAR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 115
box 378 115 478 153
use SUNSAR_cut_M1M4_2x1 xcut3 
transform 1 0 378 0 1 27
box 378 27 478 65
<< labels >>
flabel m3 s 774 0 874 176 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m3 s 378 0 478 176 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
