magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 3636 480
<< m1 >>
rect 54 -20 3618 20
rect 3582 20 3618 60
rect 54 60 3546 100
rect 3582 60 3618 100
rect 54 100 90 140
rect 3582 100 3618 140
rect 54 140 90 180
rect 126 140 3618 180
rect 54 180 90 220
rect 3582 180 3618 220
rect 54 220 3546 260
rect 3582 220 3618 260
rect 54 260 90 300
rect 3582 260 3618 300
rect 54 300 90 340
rect 126 300 3618 340
rect 54 340 90 380
rect 54 380 3618 420
<< m2 >>
rect 54 -20 3618 20
rect 3582 20 3618 60
rect 54 60 3546 100
rect 3582 60 3618 100
rect 54 100 90 140
rect 3582 100 3618 140
rect 54 140 90 180
rect 126 140 3618 180
rect 54 180 90 220
rect 3582 180 3618 220
rect 54 220 3546 260
rect 3582 220 3618 260
rect 54 260 90 300
rect 3582 260 3618 300
rect 54 300 90 340
rect 126 300 3618 340
rect 54 340 90 380
rect 54 380 3618 420
<< locali >>
rect 54 -20 3618 20
rect 3582 20 3618 60
rect 54 60 3546 100
rect 3582 60 3618 100
rect 54 100 90 140
rect 3582 100 3618 140
rect 54 140 90 180
rect 126 140 3618 180
rect 54 180 90 220
rect 3582 180 3618 220
rect 54 220 3546 260
rect 3582 220 3618 260
rect 54 260 90 300
rect 3582 260 3618 300
rect 54 300 90 340
rect 126 300 3618 340
rect 54 340 90 380
rect 54 380 3618 420
<< v1 >>
rect 3438 -16 3474 -12
rect 3438 -12 3474 -8
rect 3438 -8 3474 -4
rect 3438 -4 3474 0
rect 3438 0 3474 4
rect 3438 4 3474 8
rect 3438 8 3474 12
rect 3438 12 3474 16
rect 3474 -16 3510 -12
rect 3474 -12 3510 -8
rect 3474 -8 3510 -4
rect 3474 -4 3510 0
rect 3474 0 3510 4
rect 3474 4 3510 8
rect 3474 8 3510 12
rect 3474 12 3510 16
rect 3510 -16 3546 -12
rect 3510 -12 3546 -8
rect 3510 -8 3546 -4
rect 3510 -4 3546 0
rect 3510 0 3546 4
rect 3510 4 3546 8
rect 3510 8 3546 12
rect 3510 12 3546 16
rect 162 64 198 68
rect 162 68 198 72
rect 162 72 198 76
rect 162 76 198 80
rect 162 80 198 84
rect 162 84 198 88
rect 162 88 198 92
rect 162 92 198 96
rect 198 64 234 68
rect 198 68 234 72
rect 198 72 234 76
rect 198 76 234 80
rect 198 80 234 84
rect 198 84 234 88
rect 198 88 234 92
rect 198 92 234 96
rect 234 64 270 68
rect 234 68 270 72
rect 234 72 270 76
rect 234 76 270 80
rect 234 80 270 84
rect 234 84 270 88
rect 234 88 270 92
rect 234 92 270 96
rect 3438 144 3474 148
rect 3438 148 3474 152
rect 3438 152 3474 156
rect 3438 156 3474 160
rect 3438 160 3474 164
rect 3438 164 3474 168
rect 3438 168 3474 172
rect 3438 172 3474 176
rect 3474 144 3510 148
rect 3474 148 3510 152
rect 3474 152 3510 156
rect 3474 156 3510 160
rect 3474 160 3510 164
rect 3474 164 3510 168
rect 3474 168 3510 172
rect 3474 172 3510 176
rect 3510 144 3546 148
rect 3510 148 3546 152
rect 3510 152 3546 156
rect 3510 156 3546 160
rect 3510 160 3546 164
rect 3510 164 3546 168
rect 3510 168 3546 172
rect 3510 172 3546 176
rect 162 224 198 228
rect 162 228 198 232
rect 162 232 198 236
rect 162 236 198 240
rect 162 240 198 244
rect 162 244 198 248
rect 162 248 198 252
rect 162 252 198 256
rect 198 224 234 228
rect 198 228 234 232
rect 198 232 234 236
rect 198 236 234 240
rect 198 240 234 244
rect 198 244 234 248
rect 198 248 234 252
rect 198 252 234 256
rect 234 224 270 228
rect 234 228 270 232
rect 234 232 270 236
rect 234 236 270 240
rect 234 240 270 244
rect 234 244 270 248
rect 234 248 270 252
rect 234 252 270 256
rect 3438 304 3474 308
rect 3438 308 3474 312
rect 3438 312 3474 316
rect 3438 316 3474 320
rect 3438 320 3474 324
rect 3438 324 3474 328
rect 3438 328 3474 332
rect 3438 332 3474 336
rect 3474 304 3510 308
rect 3474 308 3510 312
rect 3474 312 3510 316
rect 3474 316 3510 320
rect 3474 320 3510 324
rect 3474 324 3510 328
rect 3474 328 3510 332
rect 3474 332 3510 336
rect 3510 304 3546 308
rect 3510 308 3546 312
rect 3510 312 3546 316
rect 3510 316 3546 320
rect 3510 320 3546 324
rect 3510 324 3546 328
rect 3510 328 3546 332
rect 3510 332 3546 336
rect 162 384 198 388
rect 162 388 198 392
rect 162 392 198 396
rect 162 396 198 400
rect 162 400 198 404
rect 162 404 198 408
rect 162 408 198 412
rect 162 412 198 416
rect 198 384 234 388
rect 198 388 234 392
rect 198 392 234 396
rect 198 396 234 400
rect 198 400 234 404
rect 198 404 234 408
rect 198 408 234 412
rect 198 412 234 416
rect 234 384 270 388
rect 234 388 270 392
rect 234 392 270 396
rect 234 396 270 400
rect 234 400 270 404
rect 234 404 270 408
rect 234 408 270 412
rect 234 412 270 416
<< v2 >>
rect 3438 -16 3474 -12
rect 3438 -12 3474 -8
rect 3438 -8 3474 -4
rect 3438 -4 3474 0
rect 3438 0 3474 4
rect 3438 4 3474 8
rect 3438 8 3474 12
rect 3438 12 3474 16
rect 3474 -16 3510 -12
rect 3474 -12 3510 -8
rect 3474 -8 3510 -4
rect 3474 -4 3510 0
rect 3474 0 3510 4
rect 3474 4 3510 8
rect 3474 8 3510 12
rect 3474 12 3510 16
rect 3510 -16 3546 -12
rect 3510 -12 3546 -8
rect 3510 -8 3546 -4
rect 3510 -4 3546 0
rect 3510 0 3546 4
rect 3510 4 3546 8
rect 3510 8 3546 12
rect 3510 12 3546 16
rect 162 64 198 68
rect 162 68 198 72
rect 162 72 198 76
rect 162 76 198 80
rect 162 80 198 84
rect 162 84 198 88
rect 162 88 198 92
rect 162 92 198 96
rect 198 64 234 68
rect 198 68 234 72
rect 198 72 234 76
rect 198 76 234 80
rect 198 80 234 84
rect 198 84 234 88
rect 198 88 234 92
rect 198 92 234 96
rect 234 64 270 68
rect 234 68 270 72
rect 234 72 270 76
rect 234 76 270 80
rect 234 80 270 84
rect 234 84 270 88
rect 234 88 270 92
rect 234 92 270 96
rect 3438 144 3474 148
rect 3438 148 3474 152
rect 3438 152 3474 156
rect 3438 156 3474 160
rect 3438 160 3474 164
rect 3438 164 3474 168
rect 3438 168 3474 172
rect 3438 172 3474 176
rect 3474 144 3510 148
rect 3474 148 3510 152
rect 3474 152 3510 156
rect 3474 156 3510 160
rect 3474 160 3510 164
rect 3474 164 3510 168
rect 3474 168 3510 172
rect 3474 172 3510 176
rect 3510 144 3546 148
rect 3510 148 3546 152
rect 3510 152 3546 156
rect 3510 156 3546 160
rect 3510 160 3546 164
rect 3510 164 3546 168
rect 3510 168 3546 172
rect 3510 172 3546 176
rect 162 224 198 228
rect 162 228 198 232
rect 162 232 198 236
rect 162 236 198 240
rect 162 240 198 244
rect 162 244 198 248
rect 162 248 198 252
rect 162 252 198 256
rect 198 224 234 228
rect 198 228 234 232
rect 198 232 234 236
rect 198 236 234 240
rect 198 240 234 244
rect 198 244 234 248
rect 198 248 234 252
rect 198 252 234 256
rect 234 224 270 228
rect 234 228 270 232
rect 234 232 270 236
rect 234 236 270 240
rect 234 240 270 244
rect 234 244 270 248
rect 234 248 270 252
rect 234 252 270 256
rect 3438 304 3474 308
rect 3438 308 3474 312
rect 3438 312 3474 316
rect 3438 316 3474 320
rect 3438 320 3474 324
rect 3438 324 3474 328
rect 3438 328 3474 332
rect 3438 332 3474 336
rect 3474 304 3510 308
rect 3474 308 3510 312
rect 3474 312 3510 316
rect 3474 316 3510 320
rect 3474 320 3510 324
rect 3474 324 3510 328
rect 3474 328 3510 332
rect 3474 332 3510 336
rect 3510 304 3546 308
rect 3510 308 3546 312
rect 3510 312 3546 316
rect 3510 316 3546 320
rect 3510 320 3546 324
rect 3510 324 3546 328
rect 3510 328 3546 332
rect 3510 332 3546 336
rect 162 384 198 388
rect 162 388 198 392
rect 162 392 198 396
rect 162 396 198 400
rect 162 400 198 404
rect 162 404 198 408
rect 162 408 198 412
rect 162 412 198 416
rect 198 384 234 388
rect 198 388 234 392
rect 198 392 234 396
rect 198 396 234 400
rect 198 400 234 404
rect 198 404 234 408
rect 198 408 234 412
rect 198 412 234 416
rect 234 384 270 388
rect 234 388 270 392
rect 234 392 270 396
rect 234 396 270 400
rect 234 400 270 404
rect 234 404 270 408
rect 234 408 270 412
rect 234 412 270 416
<< viali >>
rect 3438 -16 3474 -12
rect 3438 -12 3474 -8
rect 3438 -8 3474 -4
rect 3438 -4 3474 0
rect 3438 0 3474 4
rect 3438 4 3474 8
rect 3438 8 3474 12
rect 3438 12 3474 16
rect 3474 -16 3510 -12
rect 3474 -12 3510 -8
rect 3474 -8 3510 -4
rect 3474 -4 3510 0
rect 3474 0 3510 4
rect 3474 4 3510 8
rect 3474 8 3510 12
rect 3474 12 3510 16
rect 3510 -16 3546 -12
rect 3510 -12 3546 -8
rect 3510 -8 3546 -4
rect 3510 -4 3546 0
rect 3510 0 3546 4
rect 3510 4 3546 8
rect 3510 8 3546 12
rect 3510 12 3546 16
rect 162 64 198 68
rect 162 68 198 72
rect 162 72 198 76
rect 162 76 198 80
rect 162 80 198 84
rect 162 84 198 88
rect 162 88 198 92
rect 162 92 198 96
rect 198 64 234 68
rect 198 68 234 72
rect 198 72 234 76
rect 198 76 234 80
rect 198 80 234 84
rect 198 84 234 88
rect 198 88 234 92
rect 198 92 234 96
rect 234 64 270 68
rect 234 68 270 72
rect 234 72 270 76
rect 234 76 270 80
rect 234 80 270 84
rect 234 84 270 88
rect 234 88 270 92
rect 234 92 270 96
rect 3438 144 3474 148
rect 3438 148 3474 152
rect 3438 152 3474 156
rect 3438 156 3474 160
rect 3438 160 3474 164
rect 3438 164 3474 168
rect 3438 168 3474 172
rect 3438 172 3474 176
rect 3474 144 3510 148
rect 3474 148 3510 152
rect 3474 152 3510 156
rect 3474 156 3510 160
rect 3474 160 3510 164
rect 3474 164 3510 168
rect 3474 168 3510 172
rect 3474 172 3510 176
rect 3510 144 3546 148
rect 3510 148 3546 152
rect 3510 152 3546 156
rect 3510 156 3546 160
rect 3510 160 3546 164
rect 3510 164 3546 168
rect 3510 168 3546 172
rect 3510 172 3546 176
rect 162 224 198 228
rect 162 228 198 232
rect 162 232 198 236
rect 162 236 198 240
rect 162 240 198 244
rect 162 244 198 248
rect 162 248 198 252
rect 162 252 198 256
rect 198 224 234 228
rect 198 228 234 232
rect 198 232 234 236
rect 198 236 234 240
rect 198 240 234 244
rect 198 244 234 248
rect 198 248 234 252
rect 198 252 234 256
rect 234 224 270 228
rect 234 228 270 232
rect 234 232 270 236
rect 234 236 270 240
rect 234 240 270 244
rect 234 244 270 248
rect 234 248 270 252
rect 234 252 270 256
rect 3438 304 3474 308
rect 3438 308 3474 312
rect 3438 312 3474 316
rect 3438 316 3474 320
rect 3438 320 3474 324
rect 3438 324 3474 328
rect 3438 328 3474 332
rect 3438 332 3474 336
rect 3474 304 3510 308
rect 3474 308 3510 312
rect 3474 312 3510 316
rect 3474 316 3510 320
rect 3474 320 3510 324
rect 3474 324 3510 328
rect 3474 328 3510 332
rect 3474 332 3510 336
rect 3510 304 3546 308
rect 3510 308 3546 312
rect 3510 312 3546 316
rect 3510 316 3546 320
rect 3510 320 3546 324
rect 3510 324 3546 328
rect 3510 328 3546 332
rect 3510 332 3546 336
rect 162 384 198 388
rect 162 388 198 392
rect 162 392 198 396
rect 162 396 198 400
rect 162 400 198 404
rect 162 404 198 408
rect 162 408 198 412
rect 162 412 198 416
rect 198 384 234 388
rect 198 388 234 392
rect 198 392 234 396
rect 198 396 234 400
rect 198 400 234 404
rect 198 404 234 408
rect 198 408 234 412
rect 198 412 234 416
rect 234 384 270 388
rect 234 388 270 392
rect 234 392 270 396
rect 234 396 270 400
rect 234 400 270 404
rect 234 404 270 408
rect 234 408 270 412
rect 234 412 270 416
<< m3 >>
rect 54 -20 3618 20
rect 54 -20 3618 20
rect 3582 20 3618 60
rect 54 60 3438 100
rect 3474 60 3546 100
rect 3582 60 3618 100
rect 54 100 90 140
rect 3582 100 3618 140
rect 54 140 90 180
rect 126 140 162 180
rect 198 140 3618 180
rect 54 180 90 220
rect 3582 180 3618 220
rect 54 220 3546 260
rect 3582 220 3618 260
rect 54 260 90 300
rect 3582 260 3618 300
rect 54 300 90 340
rect 126 300 3618 340
rect 54 340 90 380
rect 54 380 3618 420
rect 54 380 3618 420
<< rm3 >>
rect 3438 60 3474 100
rect 162 140 198 180
<< v3 >>
rect 3438 -16 3474 -12
rect 3438 -12 3474 -8
rect 3438 -8 3474 -4
rect 3438 -4 3474 0
rect 3438 0 3474 4
rect 3438 4 3474 8
rect 3438 8 3474 12
rect 3438 12 3474 16
rect 3474 -16 3510 -12
rect 3474 -12 3510 -8
rect 3474 -8 3510 -4
rect 3474 -4 3510 0
rect 3474 0 3510 4
rect 3474 4 3510 8
rect 3474 8 3510 12
rect 3474 12 3510 16
rect 3510 -16 3546 -12
rect 3510 -12 3546 -8
rect 3510 -8 3546 -4
rect 3510 -4 3546 0
rect 3510 0 3546 4
rect 3510 4 3546 8
rect 3510 8 3546 12
rect 3510 12 3546 16
rect 162 64 198 68
rect 162 68 198 72
rect 162 72 198 76
rect 162 76 198 80
rect 162 80 198 84
rect 162 84 198 88
rect 162 88 198 92
rect 162 92 198 96
rect 198 64 234 68
rect 198 68 234 72
rect 198 72 234 76
rect 198 76 234 80
rect 198 80 234 84
rect 198 84 234 88
rect 198 88 234 92
rect 198 92 234 96
rect 234 64 270 68
rect 234 68 270 72
rect 234 72 270 76
rect 234 76 270 80
rect 234 80 270 84
rect 234 84 270 88
rect 234 88 270 92
rect 234 92 270 96
rect 3438 144 3474 148
rect 3438 148 3474 152
rect 3438 152 3474 156
rect 3438 156 3474 160
rect 3438 160 3474 164
rect 3438 164 3474 168
rect 3438 168 3474 172
rect 3438 172 3474 176
rect 3474 144 3510 148
rect 3474 148 3510 152
rect 3474 152 3510 156
rect 3474 156 3510 160
rect 3474 160 3510 164
rect 3474 164 3510 168
rect 3474 168 3510 172
rect 3474 172 3510 176
rect 3510 144 3546 148
rect 3510 148 3546 152
rect 3510 152 3546 156
rect 3510 156 3546 160
rect 3510 160 3546 164
rect 3510 164 3546 168
rect 3510 168 3546 172
rect 3510 172 3546 176
rect 162 224 198 228
rect 162 228 198 232
rect 162 232 198 236
rect 162 236 198 240
rect 162 240 198 244
rect 162 244 198 248
rect 162 248 198 252
rect 162 252 198 256
rect 198 224 234 228
rect 198 228 234 232
rect 198 232 234 236
rect 198 236 234 240
rect 198 240 234 244
rect 198 244 234 248
rect 198 248 234 252
rect 198 252 234 256
rect 234 224 270 228
rect 234 228 270 232
rect 234 232 270 236
rect 234 236 270 240
rect 234 240 270 244
rect 234 244 270 248
rect 234 248 270 252
rect 234 252 270 256
rect 3438 304 3474 308
rect 3438 308 3474 312
rect 3438 312 3474 316
rect 3438 316 3474 320
rect 3438 320 3474 324
rect 3438 324 3474 328
rect 3438 328 3474 332
rect 3438 332 3474 336
rect 3474 304 3510 308
rect 3474 308 3510 312
rect 3474 312 3510 316
rect 3474 316 3510 320
rect 3474 320 3510 324
rect 3474 324 3510 328
rect 3474 328 3510 332
rect 3474 332 3510 336
rect 3510 304 3546 308
rect 3510 308 3546 312
rect 3510 312 3546 316
rect 3510 316 3546 320
rect 3510 320 3546 324
rect 3510 324 3546 328
rect 3510 328 3546 332
rect 3510 332 3546 336
rect 162 384 198 388
rect 162 388 198 392
rect 162 392 198 396
rect 162 396 198 400
rect 162 400 198 404
rect 162 404 198 408
rect 162 408 198 412
rect 162 412 198 416
rect 198 384 234 388
rect 198 388 234 392
rect 198 392 234 396
rect 198 396 234 400
rect 198 400 234 404
rect 198 404 234 408
rect 198 408 234 412
rect 198 412 234 416
rect 234 384 270 388
rect 234 388 270 392
rect 234 392 270 396
rect 234 396 270 400
rect 234 400 270 404
rect 234 404 270 408
rect 234 408 270 412
rect 234 412 270 416
<< m4 >>
rect 54 -20 3618 20
rect 3582 20 3618 60
rect 54 60 3546 100
rect 3582 60 3618 100
rect 54 100 90 140
rect 3582 100 3618 140
rect 54 140 90 180
rect 126 140 3618 180
rect 54 180 90 220
rect 3582 180 3618 220
rect 54 220 3546 260
rect 3582 220 3618 260
rect 54 260 90 300
rect 3582 260 3618 300
rect 54 300 90 340
rect 126 300 3618 340
rect 54 340 90 380
rect 54 380 3618 420
<< labels >>
flabel m3 s 54 -20 3618 20 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 54 380 3618 420 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3636 480
<< end >>
