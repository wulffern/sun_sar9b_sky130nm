magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 1260 1936
<< locali >>
rect 828 291 912 325
rect 912 389 1020 423
rect 912 291 946 423
rect 990 423 1044 457
rect 828 467 912 501
rect 912 687 1044 721
rect 912 1655 1044 1689
rect 912 467 946 1689
rect 216 951 300 985
rect 300 467 432 501
rect 300 467 334 985
rect 240 1357 300 1391
rect 300 467 432 501
rect 300 467 334 1391
rect 216 1391 270 1425
rect 432 731 516 765
rect 432 995 516 1029
rect 516 731 550 1029
rect 432 1435 516 1469
rect 432 1699 516 1733
rect 516 1435 550 1733
rect 216 1831 300 1865
rect 300 1699 432 1733
rect 300 1699 334 1865
rect 162 599 270 633
rect 162 247 270 281
rect 378 1875 486 1909
rect 378 1699 486 1733
<< m1 >>
rect 1044 951 1128 985
rect 1044 1391 1128 1425
rect 828 291 1128 325
rect 1128 291 1162 1425
rect 240 653 300 687
rect 300 291 432 325
rect 300 291 334 687
rect 216 687 270 721
rect 216 1655 300 1689
rect 300 1391 1044 1425
rect 300 1391 334 1689
rect 216 1127 300 1161
rect 300 995 432 1029
rect 300 995 334 1161
rect 828 1171 912 1205
rect 912 863 1044 897
rect 912 1303 1044 1337
rect 912 863 946 1337
rect 828 1875 912 1909
rect 912 1567 1044 1601
rect 912 1567 946 1909
<< m3 >>
rect 774 0 874 1936
rect 378 0 478 1936
rect 774 0 874 1936
rect 378 0 478 1936
use SUNSAR_TAPCELLB_CV XA0 
transform 1 0 0 0 1 0
box 0 0 1260 176
use SUNSAR_IVX1_CV XA1 
transform 1 0 0 0 1 176
box 0 176 1260 352
use SUNSAR_IVX1_CV XA2 
transform 1 0 0 0 1 352
box 0 352 1260 528
use SUNSAR_IVTRIX1_CV XA3 
transform 1 0 0 0 1 528
box 0 528 1260 792
use SUNSAR_IVTRIX1_CV XA4 
transform 1 0 0 0 1 792
box 0 792 1260 1056
use SUNSAR_IVX1_CV XA5 
transform 1 0 0 0 1 1056
box 0 1056 1260 1232
use SUNSAR_IVTRIX1_CV XA6 
transform 1 0 0 0 1 1232
box 0 1232 1260 1496
use SUNSAR_IVTRIX1_CV XA7 
transform 1 0 0 0 1 1496
box 0 1496 1260 1760
use SUNSAR_IVX1_CV XA8 
transform 1 0 0 0 1 1760
box 0 1760 1260 1936
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 990 0 1 951
box 990 951 1082 985
use SUNSAR_cut_M1M2_2x1 xcut1 
transform 1 0 990 0 1 1391
box 990 1391 1082 1425
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 774 0 1 291
box 774 291 866 325
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 162 0 1 687
box 162 687 254 721
use SUNSAR_cut_M1M2_2x1 xcut4 
transform 1 0 378 0 1 291
box 378 291 470 325
use SUNSAR_cut_M1M2_2x1 xcut5 
transform 1 0 162 0 1 1655
box 162 1655 254 1689
use SUNSAR_cut_M1M2_2x1 xcut6 
transform 1 0 990 0 1 1391
box 990 1391 1082 1425
use SUNSAR_cut_M1M2_2x1 xcut7 
transform 1 0 162 0 1 1127
box 162 1127 254 1161
use SUNSAR_cut_M1M2_2x1 xcut8 
transform 1 0 378 0 1 995
box 378 995 470 1029
use SUNSAR_cut_M1M2_2x1 xcut9 
transform 1 0 774 0 1 1171
box 774 1171 866 1205
use SUNSAR_cut_M1M2_2x1 xcut10 
transform 1 0 990 0 1 863
box 990 863 1082 897
use SUNSAR_cut_M1M2_2x1 xcut11 
transform 1 0 990 0 1 1303
box 990 1303 1082 1337
use SUNSAR_cut_M1M2_2x1 xcut12 
transform 1 0 774 0 1 1875
box 774 1875 866 1909
use SUNSAR_cut_M1M2_2x1 xcut13 
transform 1 0 990 0 1 1567
box 990 1567 1082 1601
<< labels >>
flabel locali s 162 599 270 633 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 378 1875 486 1909 0 FreeSans 400 0 0 0 Q
port 3 nsew signal bidirectional
flabel locali s 378 1699 486 1733 0 FreeSans 400 0 0 0 QN
port 4 nsew signal bidirectional
flabel m3 s 774 0 874 1936 0 FreeSans 400 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel m3 s 378 0 478 1936 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 1936
<< end >>
