magic
tech sky130A
magscale 1 1
timestamp 1712786400
<< checkpaint >>
rect 0 0 1260 1760
<< locali >>
rect 1044 247 1128 281
rect 1044 1303 1128 1337
rect 1044 1655 1128 1689
rect 1128 247 1162 1689
rect 240 917 300 951
rect 300 819 432 853
rect 300 819 334 951
rect 236 951 270 985
rect 216 1567 300 1601
rect 300 995 432 1029
rect 300 995 334 1601
rect 216 1215 300 1249
rect 300 995 432 1029
rect 300 995 334 1249
rect 98 423 216 457
rect 98 1479 216 1513
rect 98 423 132 1513
rect 162 1127 270 1161
rect 990 1655 1098 1689
rect 162 247 270 281
rect 162 1479 270 1513
rect 378 1347 486 1381
rect 378 1699 486 1733
rect 774 379 882 413
<< m1 >>
rect 216 599 300 633
rect 216 1127 300 1161
rect 300 599 334 1161
rect 98 247 216 281
rect 98 1655 216 1689
rect 98 1303 216 1337
rect 98 247 132 1689
<< m3 >>
rect 774 0 866 1760
rect 378 0 470 1760
rect 774 0 866 1760
rect 378 0 470 1760
use SUNSAR_TAPCELLB_CV XA0 
transform 1 0 0 0 1 0
box 0 0 1260 176
use SUNSAR_SAREMX1_CV XA1 
transform 1 0 0 0 1 176
box 0 176 1260 880
use SUNSAR_IVX1_CV XA2 
transform 1 0 0 0 1 880
box 0 880 1260 1056
use SUNSAR_SARLTX1_CV XA4 
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNSAR_SARLTX1_CV XA5 
transform 1 0 0 0 1 1408
box 0 1408 1260 1760
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 178 0 1 599
box 178 599 270 633
use SUNSAR_cut_M1M2_2x1 xcut1 
transform 1 0 178 0 1 1127
box 178 1127 270 1161
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 162 0 1 247
box 162 247 254 281
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 162 0 1 1655
box 162 1655 254 1689
use SUNSAR_cut_M1M2_2x1 xcut4 
transform 1 0 162 0 1 1303
box 162 1303 254 1337
<< labels >>
flabel locali s 162 1127 270 1161 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew signal bidirectional
flabel locali s 990 1655 1098 1689 0 FreeSans 400 0 0 0 RST_N
port 4 nsew signal bidirectional
flabel locali s 162 247 270 281 0 FreeSans 400 0 0 0 EN
port 3 nsew signal bidirectional
flabel locali s 162 1479 270 1513 0 FreeSans 400 0 0 0 CMP_ON
port 2 nsew signal bidirectional
flabel locali s 378 1347 486 1381 0 FreeSans 400 0 0 0 CHL_OP
port 6 nsew signal bidirectional
flabel locali s 378 1699 486 1733 0 FreeSans 400 0 0 0 CHL_ON
port 7 nsew signal bidirectional
flabel locali s 774 379 882 413 0 FreeSans 400 0 0 0 ENO
port 5 nsew signal bidirectional
flabel m3 s 774 0 866 1760 0 FreeSans 400 0 0 0 AVDD
port 8 nsew signal bidirectional
flabel m3 s 378 0 470 1760 0 FreeSans 400 0 0 0 AVSS
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 1760
<< end >>
