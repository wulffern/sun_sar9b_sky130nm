magic
tech sky130A
magscale 1 1
timestamp 1712959200
<< checkpaint >>
rect 0 0 34 92
<< locali >>
rect 0 0 34 92
<< viali >>
rect 3 6 31 34
rect 3 58 31 86
<< m1 >>
rect 0 0 34 92
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 34 92
<< end >>
