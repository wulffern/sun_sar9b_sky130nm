magic
tech sky130A
magscale 1 2
timestamp 1713029161
<< locali >>
rect 168 3124 1440 3192
rect 168 2664 236 3124
rect 628 2694 864 2762
rect 0 2596 236 2664
rect 398 1550 466 2674
rect 628 2410 696 2694
rect 756 2518 1100 2586
rect 628 2342 864 2410
rect 628 2058 696 2342
rect 1032 2234 1100 2518
rect 864 2166 1100 2234
rect 628 1990 864 2058
rect 628 1706 696 1990
rect 1032 1882 1100 2166
rect 864 1814 1100 1882
rect 628 1638 864 1706
rect 628 1354 696 1638
rect 1032 1530 1100 1814
rect 864 1462 1100 1530
rect 628 1286 864 1354
rect 398 142 466 1266
rect 628 1002 696 1286
rect 756 1110 1100 1178
rect 628 934 864 1002
rect 628 650 696 934
rect 1032 826 1100 1110
rect 3420 846 3636 914
rect 864 758 1100 826
rect 628 582 864 650
rect 628 298 696 582
rect 1032 474 1100 758
rect 1764 494 1980 562
rect 864 406 1100 474
rect 628 230 864 298
rect 1032 122 1100 406
rect 864 54 1100 122
<< metal1 >>
rect 600 2870 2304 2938
rect 600 2674 668 2870
rect 432 2606 668 2674
rect 2040 2200 3096 2268
rect 2040 1794 2108 2200
rect 1872 1726 2108 1794
rect 2988 1638 3420 1706
rect 1032 1286 2304 1354
rect 1032 1002 1100 1286
rect 864 934 1100 1002
rect 3264 846 3528 914
rect 3264 650 3332 846
rect 3096 582 3332 650
<< metal2 >>
rect 1432 1814 2304 1882
rect 1432 914 1500 1814
rect 1872 1550 2108 1618
rect 432 846 1500 914
rect 2040 684 2108 1550
rect 3096 1110 3332 1178
rect 2040 616 2304 684
rect 3264 28 3332 1110
rect 3264 -40 4376 28
<< metal3 >>
rect 1676 2870 1860 2938
rect 788 230 972 298
rect 2196 0 2380 4800
rect 2988 0 3172 4800
rect 4156 2680 7848 2748
rect 4156 1706 4224 2680
rect 3512 1638 4224 1706
use SUNSAR_NCHDLR  M1
timestamp 1712959200
transform 1 0 0 0 1 0
box -180 -132 1260 484
use SUNSAR_NCHDLR  M2
timestamp 1712959200
transform 1 0 0 0 1 352
box -180 -132 1260 484
use SUNSAR_NCHDLR  M3
timestamp 1712959200
transform 1 0 0 0 1 704
box -180 -132 1260 484
use SUNSAR_NCHDLR  M4
timestamp 1712959200
transform 1 0 0 0 1 1056
box -180 -132 1260 484
use SUNSAR_NCHDLR  M5
timestamp 1712959200
transform 1 0 0 0 1 1408
box -180 -132 1260 484
use SUNSAR_NCHDLR  M6
timestamp 1712959200
transform 1 0 0 0 1 1760
box -180 -132 1260 484
use SUNSAR_NCHDLR  M7
timestamp 1712959200
transform 1 0 0 0 1 2112
box -180 -132 1260 484
use SUNSAR_NCHDLR  M8
timestamp 1712959200
transform 1 0 0 0 1 2464
box -180 -132 1260 484
use SUNSAR_IVX1_CV  XA0
timestamp 1713029161
transform 1 0 1440 0 1 352
box -180 -132 2700 484
use SUNSAR_TIEH_CV  XA1
timestamp 1713029161
transform 1 0 1440 0 1 1936
box -180 -132 2700 484
use SUNSAR_TIEL_CV  XA2
timestamp 1713029161
transform 1 0 1440 0 1 2640
box -180 -132 2700 484
use SUNSAR_TGPD_CV  XA3
timestamp 1713029161
transform 1 0 1440 0 1 704
box -180 -132 2700 836
use SUNSAR_SARBSSWCTRL_CV  XA4
timestamp 1713029161
transform 1 0 1440 0 1 1408
box -180 -132 2700 660
use SUNSAR_TAPCELLB_CV  XA5
timestamp 1713029161
transform 1 0 1440 0 1 2992
box -180 -132 2700 484
use SUNSAR_TAPCELLB_CV  XA5b
timestamp 1713029161
transform 1 0 1440 0 1 0
box -180 -132 2700 484
use SUNSAR_TAPCELLB_CV  XA7
timestamp 1713029161
transform 1 0 1440 0 1 2288
box -180 -132 2700 484
use SUNSAR_CAP_BSSW5_CV  XCAPB1
timestamp 1713029161
transform 1 0 4176 0 1 0
box -20 -51 7364 4691
use SUNSAR_cut_M1M2_2x1  xcut0
timestamp 1712959200
transform 1 0 2988 0 1 1638
box 0 0 184 68
use SUNSAR_cut_M2M4_2x1  xcut1
timestamp 1712959200
transform 1 0 3420 0 1 1638
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut2
timestamp 1712959200
transform 1 0 2988 0 1 582
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut3
timestamp 1712959200
transform 1 0 3420 0 1 846
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut4
timestamp 1712959200
transform 1 0 1764 0 1 1550
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut5
timestamp 1712959200
transform 1 0 2196 0 1 616
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut6
timestamp 1712959200
transform 1 0 324 0 1 2606
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut7
timestamp 1712959200
transform 1 0 2196 0 1 2870
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut8
timestamp 1712959200
transform 1 0 1764 0 1 1726
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut9
timestamp 1712959200
transform 1 0 2988 0 1 2200
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut10
timestamp 1712959200
transform 1 0 756 0 1 934
box 0 0 184 68
use SUNSAR_cut_M1M2_2x1  xcut11
timestamp 1712959200
transform 1 0 2196 0 1 1286
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut12
timestamp 1712959200
transform 1 0 2228 0 1 1814
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut13
timestamp 1712959200
transform 1 0 356 0 1 846
box 0 0 184 68
use SUNSAR_cut_M1M3_2x1  xcut14
timestamp 1712959200
transform 1 0 2988 0 1 1110
box 0 0 184 68
use SUNSAR_cut_M3M4_2x1  xcut15
timestamp 1712959200
transform 1 0 4284 0 1 -40
box 0 0 184 68
use SUNSAR_cut_M1M4_2x1  xcut16
timestamp 1712959200
transform 1 0 788 0 1 230
box 0 0 184 68
use SUNSAR_cut_M2M4_2x1  xcut17
timestamp 1712959200
transform 1 0 1676 0 1 2870
box 0 0 184 68
<< labels >>
flabel metal3 s 788 230 972 298 0 FreeSans 800 0 0 0 VI
port 1 nsew signal bidirectional
flabel metal3 s 1676 2870 1860 2938 0 FreeSans 800 0 0 0 TIE_L
port 4 nsew signal bidirectional
flabel locali s 1764 494 1980 562 0 FreeSans 800 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 3420 846 3636 914 0 FreeSans 800 0 0 0 CKN
port 3 nsew signal bidirectional
flabel locali s 756 1110 972 1178 0 FreeSans 800 0 0 0 VO1
port 5 nsew signal bidirectional
flabel locali s 756 2518 972 2586 0 FreeSans 800 0 0 0 VO2
port 6 nsew signal bidirectional
flabel metal3 s 2988 0 3172 4800 0 FreeSans 800 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel metal3 s 2196 0 2380 4800 0 FreeSans 800 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 11448 4800
<< end >>
