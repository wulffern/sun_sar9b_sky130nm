*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SUNSAR_SARBSSW_CV_lpe.spi
#else
.include ../../../work/xsch/SUNSAR_SARBSSW_CV.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-4

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------

.param TRF = 10p

*- Analog parameters
.param AVDD = {vdda}

*- 8 MHz clock frequency
.param PERIOD_CLK = 125n

*- 25% duty-cycle clock
.param PW_CLK = PERIOD_CLK/4

*- Frequency bin of the input signal
.param fbin = 5

*- number of cycles in FFT
.param nbpt = 128

*- Sampling frequency
.param fs = 1/PERIOD_CLK

*- Input frequency for coherent sampling
.param fin = fbin/nbpt*fs

.param vamp = 0.5

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0     dc 0
VDD  AVDD  0  pwl 0 0 10n {AVDD}

VCLK CK 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})

VCM VCM 0 dc {AVDD/2}
VSARP SAR_IP VCM sin (0 {vamp} {fin} )
VSARN SAR_IN VCM sin (0 {-vamp} {fin} )


XDUT1 SAR_IP CK CKN1 TIE_L1 SARP SARN AVDD AVSS  SUNSAR_SARBSSW_CV
XDUT2 SAR_IN CK CKN2 TIE_L1 SARN SARP AVDD AVSS  SUNSAR_SARBSSW_CV

C1 SARP 0 300f
C2 SARN 0 300f

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(SARP)
.save v(SARN)
.save v(SAR_IP)
.save v(SAR_IN)
.save v(ck)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 10n 500n 125n

let sar_in = v(sar_ip)-v(sar_in)
let sar_diff = v(sarp)-v(sarn)
let sar_cm = (v(sarp)+v(sarn))/2
write
quit


.endc

.end
