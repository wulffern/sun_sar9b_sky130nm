* NGSPICE file created from SUNSAR_SAR9B_CV.ext - technology: sky130B

.subckt SUNSAR_SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4>
+ D<3> D<2> D<1> D<0> EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
R0 XDAC1.XC128a<1>.XRES16.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X0 XB1.XA0.MP0.D CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X1 AVDD XA4.XA1.XA1.MN0.S XA4.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X2 AVSS XA8.XA3.MN0.G D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X3 XA5.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA6.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X4 XA1.XA10.MP0.G XA1.XA9.MN1.G XA1.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X5 XA0.XA12.MP0.D XA0.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X6 AVDD XA1.XA9.MN1.G XA1.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X7 VREF XA6.XA4.MN0.D XA6.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X8 VREF XA4.XA4.MN0.G XA4.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X9 XA2.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R1 XDAC1.XC64b<1>.XRES1B.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X10 XA5.XA10.MP0.D XA5.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X11 AVSS CK_SAMPLE XA1.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X12 VREF XA6.XA4.MN0.G XA6.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X13 AVDD XA1.XA6.MP0.G XA1.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X14 VREF XA4.XA3.MN0.G D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X15 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X16 XA8.XA9.MN1.G CK_SAMPLE XA8.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X17 XA5.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R2 XA0.XA6.MP0.G XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X18 VREF XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X19 XA20.XA2.MN1.D SARP XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X20 XA20.XA3a.MN0.G XA20.XA3.MN6.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X21 XA6.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X22 XA4.XA9.MN1.G D<4> XA4.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X23 AVSS XA2.XA4.MN0.D XA2.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R3 XDAC1.XC128b<2>.XRES1B.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X24 XA8.XA11.MN1.G XA7.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X25 XA5.XA10.MP0.G XA5.XA9.MN1.G XA5.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X26 XA5.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA5.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X27 XA8.XA11.MN1.G XA7.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X28 XA6.XA4.MN0.D XA6.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X29 AVDD XA20.XA9.MP0.D XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X30 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=227 pd=1.22k as=0.616 ps=3.3 w=1.08 l=0.18
X31 AVSS XA2.XA4.MN0.G XA2.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R4 XDAC1.XC32a<0>.XRES16.B D<6> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X32 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=150 pd=802 as=0.616 ps=3.3 w=1.08 l=0.18
X33 AVSS XA8.XA11.MN1.G XA8.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X34 AVSS CK_SAMPLE XA5.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X35 AVSS XA20.XA3.MN6.D XA20.XA2a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X36 AVDD XA20.XA3.MN6.D XA20.XA2a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X37 VREF XA0.XA1.XA5.MN2.D D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X38 XA20.XA1.MN0.D XA20.XA10.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X39 XA0.XA9.MN0.D XA0.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X40 AVSS XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R5 XDAC1.X16ab.XRES1B.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X41 AVDD XA20.XA10.MN1.D XA20.XA1.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R6 D<8> XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X42 XA8.XA4.MN0.G EN XA8.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X43 XA8.XA7.MP0.D XA8.XA7.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X44 XA20.XA3.MN0.D SARP XA20.XA2.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X45 AVDD XA20.XA3.MN6.D XA20.XA3a.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X46 XA0.XA1.XA4.MP1.D EN XA0.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X47 XA4.XA12.MP0.G XA4.XA11.MN1.G XA4.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X48 VREF XA5.XA4.MN0.D XA5.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X49 XA2.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X50 XA8.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA8.XA7.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X51 XA0.XA6.MP2.G D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X52 SARN XB2.M1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X53 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=7.39 ps=39.6 w=1.08 l=0.18
X54 XA6.XA10.MP0.D XA6.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X55 XA2.XA4.MN0.D XA2.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X56 AVDD XB1.XA0.MP0.D XB1.XA3.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X57 AVDD EN XA0.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X58 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X59 XA4.XA7.MP0.D XA5.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X60 VREF XA5.XA3.MN0.G D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X61 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X62 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X63 XA8.XA12.MP0.G XA8.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R7 XDAC1.XC1.XRES1B.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X64 D<8> XA0.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X65 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X66 XA6.XA6.MP2.D D<2> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X67 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X68 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X69 XA7.XA9.MN0.D XA7.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X70 XA7.XA10.MP0.G XA7.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X71 XA3.XA1.XA5.MN2.D XA3.XA1.XA5.MN2.G XA3.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X72 XA3.XA1.XA5.MN2.D EN XA3.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X73 XA0.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X74 XA4.XA11.MP0.D XA4.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X75 XA3.XA4.MN0.D XA3.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R8 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X76 XA3.XA1.XA2.MP0.D XA4.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X77 XA3.XA4.MN0.D XA3.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X78 XA3.XA1.XA2.MP0.D XA4.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X79 AVDD XA6.XA9.MN1.G XA6.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X80 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X81 XA2.XA10.MP0.D XA2.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X82 XA5.XA6.MP0.G XA5.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X83 XA8.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA8.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X84 D<5> XA3.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X85 D<5> XA3.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X86 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=7.39 ps=39.6 w=1.08 l=0.18
X87 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X88 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X89 AVDD XA6.XA6.MP0.G XA6.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X90 XA2.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X91 XA3.XA1.XA5.MN1.D XA3.XA1.XA2.MP0.D XA3.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X92 XA20.XA3.MN1.D SARN XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X93 XA3.XA1.XA5.MP1.D EN XA3.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X94 XA20.XA3.MN1.D XA20.XA9.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X95 XA6.XA4.MN0.G XA6.XA1.XA5.MN2.G XA6.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X96 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X97 XA6.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X98 AVDD XA3.XA1.XA1.MN0.S XA3.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X99 XA0.XA8.MP0.D XA0.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X100 VREF XA8.XA4.MN0.D XA8.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X101 XA2.XA10.MP0.G XA2.XA9.MN1.G XA2.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X102 VREF XA3.XA4.MN0.G XA3.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X103 AVSS XA3.XA4.MN0.G XA3.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X104 XA0.XA6.MP0.G XA0.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X105 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X106 VREF XA8.XA3.MN0.G D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X107 VREF XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X108 AVSS CK_SAMPLE XA2.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X109 AVSS XA3.XA3.MN0.G D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R9 XA0.XA6.MP0.G XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X110 VREF XA3.XA3.MN0.G D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X111 XB2.XA0.MP0.D CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X112 XA2.XA1.XA4.MP1.D EN XA2.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X113 XA6.XA11.MN1.G XA5.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X114 XA4.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X115 D<6> XA2.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X116 AVDD EN XA2.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X117 XA3.XA9.MN1.G CK_SAMPLE XA3.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X118 XA3.XA9.MN1.G D<5> XA3.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X119 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X120 AVSS XA20.XA2a.MN0.D XA6.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X121 XA8.XA6.MP0.G XA8.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X122 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R10 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R11 XDAC1.XC0.XRES2.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R12 D<8> XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X123 XA2.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X124 AVSS XA4.XA4.MN0.D XA4.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R13 XA2.XA6.MP0.G XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X125 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X126 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X127 AVSS XA3.XA11.MN1.G XA3.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X128 AVSS XA6.XA4.MN0.D XA6.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X129 XA3.XA12.MP0.G XA3.XA11.MN1.G XA3.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X130 AVSS XA4.XA4.MN0.G XA4.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X131 XA5.XA10.MP0.G XA5.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X132 XA1.XA1.XA5.MN2.D XA0.XA7.MP0.G XA1.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X133 XA3.XA7.MP0.D XA4.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X134 AVSS XA6.XA3.MN0.G D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X135 AVSS XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X136 XA1.XA1.XA5.MN2.D EN XA1.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X137 XA3.XA7.MP0.D XA4.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R14 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R15 XDAC1.XC64b<1>.XRES8.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X138 XA1.XA4.MN0.D XA1.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X139 XA1.XA4.MN0.D XA1.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R16 XB1.XA3.MN1.D m3_7544_1364# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X140 XA1.XA1.XA2.MP0.D XA2.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X141 XA1.XA1.XA2.MP0.D XA2.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X142 XA4.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R17 XB1.XA3.MN1.D m3_7544_4532# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R18 XB2.XA4.MP0.D m3_26048_3300# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X143 XA20.XA12.MP0.G XA8.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X144 XA2.XA8.MP0.D XA2.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X145 D<7> XA1.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X146 XA3.XA12.MP0.G XA3.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X147 XA0.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X148 XA4.XA4.MN0.D XA4.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X149 D<7> XA1.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X150 XA3.XA11.MP0.D XA3.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X151 XA2.XA6.MP0.G XA2.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X152 XA1.XA1.XA5.MN1.D XA1.XA1.XA2.MP0.D XA1.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X153 D<8> XA0.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X154 XA1.XA1.XA5.MP1.D EN XA1.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X155 XA6.XA6.MP0.G XA6.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X156 XA5.XA1.XA5.MN2.D XA5.XA1.XA5.MN2.G XA5.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X157 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X158 AVDD XA1.XA1.XA1.MN0.S XA1.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X159 XA5.XA4.MN0.D XA5.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X160 AVSS XA1.XA4.MN0.G XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R19 D<8> XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X161 XA5.XA1.XA2.MP0.D XA6.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X162 AVSS XA0.XA4.MN0.D XA0.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X163 VREF XA1.XA4.MN0.G XA1.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X164 XA4.XA10.MP0.D XA4.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X165 XA7.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X166 AVSS XA1.XA3.MN0.G D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X167 D<3> XA5.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R20 m3_16472_1364# XB2.XA3.MN1.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X168 XB1.XA4.MN0.D XB1.XA0.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X169 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X170 XA7.XA6.MP0.D XA7.XA6.MP0.G XA7.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X171 AVSS XA0.XA4.MN0.G XA0.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X172 VREF XA1.XA3.MN0.G D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R21 XDAC1.XC64b<1>.XRES1A.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R22 m3_16472_4532# XB2.XA3.MN1.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X173 XA4.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X174 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X175 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X176 XA5.XA1.XA5.MN1.D XA5.XA1.XA2.MP0.D XA5.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X177 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X178 XA8.XA10.MP0.G XA8.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X179 AVSS XA0.XA1.XA5.MN2.D D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X180 AVSS XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X181 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X182 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X183 XA1.XA9.MN1.G CK_SAMPLE XA1.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X184 XA1.XA9.MN1.G D<7> XA1.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X185 XA0.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X186 XA7.XA11.MN1.G XA6.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X187 XA4.XA10.MP0.G XA4.XA9.MN1.G XA4.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X188 AVSS XA7.XA4.MN0.D XA7.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X189 VREF XA7.XA4.MN0.D XA7.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X190 AVSS XA5.XA4.MN0.G XA5.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X191 SAR_IP XB1.XA3.MN0.S XB1.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X192 XA8.XA1.XA4.MN1.D XA8.XA1.XA2.MP0.D XA8.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X193 XA0.XA4.MN0.D XA0.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X194 VREF XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X195 AVSS XB1.XA0.MP0.D XB1.XA3.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X196 AVSS CK_SAMPLE XA4.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X197 AVSS XA7.XA4.MN0.G XA7.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X198 D<0> XA8.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R23 m3_n2104_2244# XB1.XA4.MP0.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X199 VREF XA7.XA4.MN0.G XA7.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X200 AVSS XA5.XA3.MN0.G D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X201 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X202 XA8.XA1.XA1.MN0.D XA8.XA1.XA5.MN2.G XA8.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R24 XDAC1.XC0.XRES4.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X203 XA6.XA1.XA5.MN2.D EN XA6.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X204 XA4.XA1.XA4.MP1.D EN XA4.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X205 AVSS XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X206 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X207 AVSS XA0.XA12.MP0.D XA1.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X208 VREF XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R25 XDAC1.X16ab.XRES1A.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X209 XA1.XA12.MP0.G XA0.XA12.MP0.D XA1.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X210 XA6.XA4.MN0.D XA6.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X211 D<4> XA4.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X212 XA6.XA1.XA2.MP0.D XA7.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X213 AVDD EN XA4.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X214 XA5.XA9.MN1.G CK_SAMPLE XA5.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X215 XA8.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X216 XA7.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X217 XA1.XA7.MP0.D XA2.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X218 XA7.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X219 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X220 XA0.XA10.MP0.D XA0.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X221 XA1.XA7.MP0.D XA2.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X222 D<2> XA6.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X223 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X224 XA7.XA4.MN0.D XA7.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X225 XA7.XA4.MN0.D XA7.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R26 XA6.XA6.MP0.G XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X226 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X227 XA6.XA1.XA5.MP1.D EN XA6.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X228 XA6.XA9.MN0.D XA6.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X229 XA0.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R27 XDAC1.XC1.XRES1A.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X230 XA4.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X231 XA2.XA1.XA5.MN2.D XA2.XA1.XA5.MN2.G XA2.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X232 XA1.XA12.MP0.G XA1.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X233 XA1.XA11.MP0.D XA1.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X234 AVDD XA6.XA1.XA1.MN0.S XA6.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X235 XA20.XA3.MN0.D XA20.XA9.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X236 AVDD XA20.XA9.MP0.D XA20.XA3.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X237 XA2.XA4.MN0.D XA2.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X238 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X239 XA2.XA1.XA2.MP0.D XA3.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X240 SARP XB1.M1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X241 AVSS XA5.XA11.MN1.G XA5.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R28 D<8> XDAC2.XC128a<1>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X242 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X243 XA0.XA10.MP0.G XA0.XA9.MN1.G XA0.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X244 VREF XA6.XA4.MN0.G XA6.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X245 D<6> XA2.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R29 XDAC1.XC64a<0>.XRES1A.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X246 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R30 XDAC1.XC0.XRES16.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X247 XA7.XA10.MP0.D XA7.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X248 DONE XA8.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X249 XA5.XA7.MP0.D XA6.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X250 XA7.XA10.MP0.D XA7.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X251 VREF XA6.XA3.MN0.G D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X252 XA0.XA4.MN0.G EN XA0.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X253 AVSS CK_SAMPLE XA0.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X254 XA2.XA1.XA5.MN1.D XA2.XA1.XA2.MP0.D XA2.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X255 XB2.XA1.MP0.D XB2.XA1.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X256 XA8.XA6.MP0.G XA8.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X257 XA7.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X258 XA7.XA6.MP2.D D<1> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X259 SARN XB2.M1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X260 XA0.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA0.XA7.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X261 XA4.XA8.MP0.D XA4.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X262 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X263 XA5.XA12.MP0.G XA5.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X264 XA5.XA6.MP0.D XA5.XA6.MP0.G XA5.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R31 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X265 XB2.XA1.MN0.D XB2.XA1.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X266 XA6.XA9.MN1.G D<2> XA6.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X267 XA4.XA6.MP0.G XA4.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X268 AVSS XA2.XA4.MN0.G XA2.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X269 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X270 XA7.XA10.MP0.G XA7.XA9.MN1.G XA7.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X271 AVDD XA7.XA9.MN1.G XA7.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X272 AVDD XB2.M1.G XB2.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X273 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X274 AVSS XA2.XA3.MN0.G D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X275 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X276 AVSS CK_SAMPLE XA7.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R32 XA3.XA6.MP0.G XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X277 AVDD XA7.XA6.MP0.G XA7.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R33 XA0.XA6.MP0.G XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X278 VREF XA5.XA4.MN0.D XA5.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X279 XB2.M1.G XB2.XA1.MP0.D XB2.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X280 XA6.XA12.MP0.G XA6.XA11.MN1.G XA6.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X281 XA0.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA0.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X282 XA2.XA9.MN1.G CK_SAMPLE XA2.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X283 VREF XA5.XA4.MN0.G XA5.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X284 XA20.XA3.MN0.D SARN XA20.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X285 AVDD AVDD XA20.XA3.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R34 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X286 XA6.XA7.MP0.D XA7.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R35 XDAC1.XC64a<0>.XRES1B.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X287 VREF XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X288 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X289 AVSS XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X290 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X291 VREF XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X292 XA5.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X293 VREF XA0.XA4.MN0.D XA0.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X294 XA3.XA1.XA4.MN1.D XA3.XA1.XA2.MP0.D XA3.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X295 XA6.XA11.MP0.D XA6.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X296 XA3.XA1.XA4.MP1.D EN XA3.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X297 AVSS XA2.XA11.MN1.G XA2.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X298 XA8.XA6.MP0.D XA8.XA6.MP0.G XA8.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X299 XA5.XA4.MN0.D XA5.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R36 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X300 D<5> XA3.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X301 XA3.XA1.XA1.MN0.D XA3.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X302 VREF D<8> XA0.XA6.MP2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X303 D<5> XA3.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X304 AVDD EN XA3.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X305 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X306 AVDD XB2.XA0.MP0.D XB2.XA3.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X307 XA2.XA4.MN0.G EN XA2.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X308 XA2.XA7.MP0.D XA3.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X309 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X310 XA20.XA3.MN1.D SARN XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X311 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X312 XA20.XA3.MN6.D XA20.XA9.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X313 XB2.XA0.MP0.D CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X314 XA2.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA3.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X315 XA3.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X316 XA3.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X317 XA2.XA12.MP0.G XA2.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X318 VREF XA8.XA4.MN0.D XA8.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X319 XA5.XA10.MP0.D XA5.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R37 D<8> XDAC2.XC128a<1>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X320 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X321 XA0.XA6.MP0.G XA0.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X322 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X323 VREF XA8.XA4.MN0.G XA8.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X324 XA5.XA6.MP2.D D<3> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X325 XA4.XA1.XA5.MN2.D XA4.XA1.XA5.MN2.G XA4.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X326 VREF XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R38 XB2.XA4.MP0.D m3_26048_132# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X327 XB1.XA1.MP0.D XB1.XA1.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X328 XA4.XA4.MN0.D XA4.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R39 XDAC1.XC128b<2>.XRES2.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X329 XA4.XA1.XA2.MP0.D XA5.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X330 XA2.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA2.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X331 XA8.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X332 AVDD XA5.XA9.MN1.G XA5.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X333 XA3.XA8.MP0.D XA3.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X334 XA20.XA10.MN1.D XA20.XA12.MP0.D XA20.XA10.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X335 XA3.XA8.MP0.D XA3.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X336 XA6.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X337 D<4> XA4.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X338 AVDD XA20.XA12.MP0.D XA20.XA10.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X339 XA8.XA4.MN0.D XA8.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X340 AVDD XA5.XA6.MP0.G XA5.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X341 XA3.XA6.MP0.G XA3.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X342 XA3.XA6.MP0.G XA3.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X343 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R40 XDAC1.X16ab.XRES2.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X344 XA4.XA1.XA5.MN1.D XA4.XA1.XA2.MP0.D XA4.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X345 AVDD XB1.M1.G XB1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R41 XA5.XA6.MP0.G XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X346 XA0.XA12.MP0.D XA0.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R42 XDAC1.XC128a<1>.XRES8.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X347 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X348 VREF XA2.XA4.MN0.D XA2.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R43 D<8> XDAC2.XC128a<1>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X349 AVSS XA6.XA4.MN0.D XA6.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X350 AVSS XA4.XA4.MN0.G XA4.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X351 VREF XA2.XA3.MN0.G D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R44 XDAC1.XC1.XRES2.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R45 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X352 XA8.XA10.MP0.D XA8.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X353 AVSS XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X354 XA20.XA11.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X355 AVSS XA6.XA4.MN0.G XA6.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X356 VREF XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X357 XA20.XA11.MP0.D CK_SAMPLE AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X358 AVSS XA4.XA3.MN0.G D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X359 XA8.XA6.MP2.D D<0> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X360 XA1.XA1.XA4.MN1.D XA1.XA1.XA2.MP0.D XA1.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X361 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X362 AVSS XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X363 XA0.XA1.XA5.MN2.D EN XA0.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R46 XDAC1.XC64a<0>.XRES8.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X364 XA1.XA1.XA4.MP1.D EN XA1.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X365 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X366 D<7> XA1.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X367 XA1.XA1.XA1.MN0.D XA0.XA7.MP0.G XA1.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X368 XA0.XA4.MN0.D XA0.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X369 D<7> XA1.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X370 AVDD EN XA1.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X371 XA0.XA1.XA2.MP0.D XA0.XA7.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X372 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X373 XA4.XA9.MN1.G CK_SAMPLE XA4.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X374 XA6.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X375 XA2.XA6.MP0.G XA2.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R47 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X376 AVDD XA8.XA9.MN1.G XA8.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X377 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X378 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X379 XA6.XA4.MN0.D XA6.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X380 XA0.XA6.MP2.G D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R48 XDAC1.XC32a<0>.XRES8.B D<4> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X381 XA0.XA10.MP0.G XA0.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R49 XA2.XA3.MN0.G XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X382 AVSS XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X383 XA1.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X384 AVDD XA8.XA6.MP0.G XA8.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X385 XA0.XA1.XA5.MN1.D XA0.XA1.XA2.MP0.D XA0.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X386 XA1.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X387 XA7.XA1.XA5.MN2.D XA7.XA1.XA5.MN2.G XA7.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R50 XA3.XA3.MN0.G XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X388 XA8.XA4.MN0.G XA8.XA1.XA5.MN2.G XA8.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X389 XA7.XA1.XA5.MN2.D EN XA7.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X390 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X391 XA5.XA1.XA4.MN1.D XA5.XA1.XA2.MP0.D XA5.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X392 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X393 XA0.XA7.MP0.G XA0.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X394 AVSS XA4.XA11.MN1.G XA4.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X395 XA7.XA4.MN0.D XA7.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X396 XA7.XA4.MN0.D XA7.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X397 D<3> XA5.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X398 XA8.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X399 XA7.XA1.XA2.MP0.D XA8.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X400 XA5.XA1.XA1.MN0.D XA5.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X401 XA7.XA1.XA2.MP0.D XA8.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X402 AVSS XA0.XA4.MN0.G XA0.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X403 XA4.XA4.MN0.G EN XA4.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X404 XA6.XA10.MP0.D XA6.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X405 XA4.XA7.MP0.D XA5.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X406 D<1> XA7.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R51 XA0.XA6.MP0.G XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X407 D<1> XA7.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X408 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X409 AVSS D<8> XA0.XA6.MP2.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X410 XA4.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA5.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X411 XA3.XA11.MN1.G XA2.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X412 XA6.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X413 XA7.XA1.XA5.MN1.D XA7.XA1.XA2.MP0.D XA7.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X414 XA1.XA8.MP0.D XA1.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X415 SARN XB2.M1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X416 XA5.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X417 XA7.XA1.XA5.MP1.D EN XA7.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X418 XA1.XA8.MP0.D XA1.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X419 XA4.XA12.MP0.G XA4.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X420 XA1.XA6.MP0.G XA1.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X421 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X422 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X423 XA1.XA6.MP0.G XA1.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R52 AVSS XDAC1.XC32a<0>.XRES1A.A sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X424 AVDD XA7.XA1.XA1.MN0.S XA7.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X425 XA0.XA9.MN1.G CK_SAMPLE XA0.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X426 XA6.XA10.MP0.G XA6.XA9.MN1.G XA6.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X427 AVSS XA7.XA4.MN0.G XA7.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X428 VREF XA7.XA4.MN0.G XA7.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X429 AVSS XA20.XA2a.MN0.D XA8.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R53 XDAC1.X16ab.XRES4.B D<5> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X430 AVSS CK_SAMPLE XA6.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X431 VREF XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X432 AVSS XA7.XA3.MN0.G D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X433 SARP XB1.M1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X434 VREF XA7.XA3.MN0.G D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R54 XDAC1.XC128a<1>.XRES1A.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X435 XA4.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA4.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X436 XA6.XA1.XA4.MP1.D EN XA6.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X437 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X438 XA5.XA8.MP0.D XA5.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R55 XDAC1.XC64b<1>.XRES4.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X439 AVSS XA0.XA11.MN1.G XA0.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X440 D<2> XA6.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X441 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X442 AVDD EN XA6.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X443 AVSS XA8.XA4.MN0.D XA8.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X444 XA5.XA6.MP0.G XA5.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X445 XA2.XA10.MP0.G XA2.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X446 XA7.XA9.MN1.G CK_SAMPLE XA7.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X447 XA7.XA9.MN1.G D<1> XA7.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X448 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X449 XA0.XA7.MP0.D XA0.XA7.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X450 AVSS XA8.XA3.MN0.G D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X451 AVSS XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X452 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X453 VREF XA4.XA4.MN0.D XA4.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X454 XA6.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X455 XA2.XA1.XA4.MN1.D XA2.XA1.XA2.MP0.D XA2.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R56 XDAC1.XC128b<2>.XRES4.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X456 XA0.XA12.MP0.G XA0.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X457 VREF XA4.XA3.MN0.G D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X458 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X459 D<6> XA2.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X460 XA2.XA1.XA1.MN0.D XA2.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X461 AVSS XA7.XA11.MN1.G XA7.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X462 XA7.XA12.MP0.G XA7.XA11.MN1.G XA7.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R57 XDAC1.XC32a<0>.XRES1B.B D<1> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X463 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X464 XB2.XA2.MN0.G XB2.XA2.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X465 XA8.XA6.MP0.G XA8.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X466 XA5.XA1.XA5.MN2.D EN XA5.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X467 XA7.XA7.MP0.D XA8.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X468 XA7.XA7.MP0.D XA8.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R58 D<8> XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X469 XA5.XA4.MN0.D XA5.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X470 XB2.XA3.MN1.D AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X471 XA2.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X472 XA5.XA1.XA2.MP0.D XA6.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X473 XA0.XA11.MN1.G XB2.XA2.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X474 XA6.XA8.MP0.D XA6.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X475 XA4.XA6.MP0.G XA4.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R59 XDAC1.XC128a<1>.XRES1B.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X476 D<3> XA5.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X477 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X478 XA7.XA12.MP0.G XA7.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X479 XB2.XA3.MN1.D XB2.XA0.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X480 XA7.XA11.MP0.D XA7.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X481 XA20.XA3.MN1.D SARN XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X482 XA6.XA6.MP0.G XA6.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X483 XA20.XA3.MN6.D XA20.XA3a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R60 XDAC1.XC1.XRES4.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X484 XA5.XA1.XA5.MP1.D EN XA5.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X485 XA20.XA3a.MN0.G XA20.XA3.MN6.D XA20.XA2.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X486 XA3.XA4.MN0.G XA3.XA1.XA5.MN2.G XA3.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X487 AVDD XA20.XA3.MN6.D XA20.XA3a.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X488 XA3.XA4.MN0.G EN XA3.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R61 XDAC1.XC128b<2>.XRES16.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R62 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X489 AVDD XA5.XA1.XA1.MN0.S XA5.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X490 XA0.XA6.MP0.D XA0.XA6.MP0.G XA0.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X491 XA3.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R63 XB1.XA3.MN1.D m3_7544_308# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X492 XA3.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA4.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X493 XA2.XA8.MP0.D XA2.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X494 VREF XA5.XA4.MN0.G XA5.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X495 XA20.XA12.MP0.G XA8.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X496 XA20.XA3.MN0.D SARN XA20.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X497 AVDD XA20.XA3a.MN0.G XA20.XA3.MN6.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X498 D<8> XA0.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R64 XB1.XA3.MN1.D m3_7544_3476# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X499 XA2.XA6.MP0.G XA2.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R65 XB2.XA4.MP0.D m3_26048_2244# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X500 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X501 AVSS XB2.XA0.MP0.D XB2.XA3.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X502 VREF XA5.XA3.MN0.G D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X503 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X504 XA5.XA11.MN1.G XA4.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X505 XA20.XA3a.MN0.D XA20.XA3a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X506 XA8.XA1.XA5.MN2.D EN XA8.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X507 VREF XA0.XA4.MN0.D XA0.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X508 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X509 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X510 XA8.XA4.MN0.D XA8.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X511 XA8.XA1.XA2.MP0.D XA8.XA7.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X512 XA5.XA9.MN1.G D<3> XA5.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X513 VREF XA0.XA4.MN0.G XA0.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X514 AVSS XA20.XA2a.MN0.D XA3.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X515 XA3.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA3.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X516 XA20.XA2.MN1.D SARP XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X517 D<0> XA8.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X518 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X519 XA20.XA2.MN1.D XA20.XA9.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X520 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R66 XDAC1.XC64b<1>.XRES2.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X521 AVSS XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R67 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X522 AVDD XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X523 VREF XA0.XA1.XA5.MN2.D D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R68 XA0.XA6.MP0.G XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X524 XA8.XA1.XA5.MP1.D EN XA8.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X525 XA8.XA9.MN0.D XA8.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R69 m3_16472_3476# XB2.XA3.MN1.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X526 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X527 XA0.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X528 AVSS XA3.XA4.MN0.D XA3.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X529 AVDD XA8.XA1.XA1.MN0.S XA8.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X530 XA5.XA12.MP0.G XA5.XA11.MN1.G XA5.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X531 VREF XA3.XA4.MN0.D XA3.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X532 XA20.XA12.MP0.D XA20.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X533 XA0.XA4.MN0.D XA0.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X534 XA20.XA12.MP0.D XA20.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X535 XA4.XA10.MP0.G XA4.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X536 VREF XA8.XA4.MN0.G XA8.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X537 AVSS XA3.XA3.MN0.G D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X538 XA5.XA7.MP0.D XA6.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X539 VREF XA3.XA3.MN0.G D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X540 AVDD XA20.XA9.MP0.D XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X541 AVSS XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X542 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X543 VREF XA8.XA3.MN0.G D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X544 XB1.XA2.MN0.G XB1.XA2.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X545 XA6.XA1.XA5.MN2.D XA6.XA1.XA5.MN2.G XA6.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R70 D<8> XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X546 XA20.XA4.MN0.D XA20.XA10.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X547 XA2.XA6.MP0.D XA2.XA6.MP0.G XA2.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R71 m3_n2104_1188# XB1.XA4.MP0.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X548 XA4.XA1.XA4.MN1.D XA4.XA1.XA2.MP0.D XA4.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X549 AVDD XA20.XA10.MN1.D XA20.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R72 m3_n2104_4356# XB1.XA4.MP0.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X550 XB1.XA3.MN1.D AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X551 XA5.XA11.MP0.D XA5.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X552 XA6.XA4.MN0.D XA6.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X553 AVSS DONE XA20.XA11.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X554 D<4> XA4.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R73 XA3.XA3.MN0.G XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X555 XA6.XA1.XA2.MP0.D XA7.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X556 XA20.XA11.MN0.D DONE XA20.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X557 XA0.XA10.MP0.D XA0.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X558 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X559 XA4.XA1.XA1.MN0.D XA4.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X560 XA8.XA9.MN1.G D<0> XA8.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X561 XA3.XA6.MP0.G XA3.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X562 XA1.XA4.MN0.G XA0.XA7.MP0.G XA1.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X563 XA3.XA6.MP0.G XA3.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X564 D<2> XA6.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X565 XA1.XA4.MN0.G EN XA1.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X566 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X567 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X568 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X569 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X570 XA0.XA6.MP2.D XA0.XA6.MP2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X571 XA1.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X572 XA20.XA3.MN6.D XA20.XA3a.MN0.G XA20.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X573 XA1.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA2.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X574 XA4.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X575 XA6.XA1.XA5.MN1.D XA6.XA1.XA2.MP0.D XA6.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X576 AVDD XA20.XA3a.MN0.G XA20.XA3.MN6.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X577 VREF XA2.XA4.MN0.D XA2.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X578 AVDD XA0.XA9.MN1.G XA0.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X579 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X580 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X581 VREF XA2.XA4.MN0.G XA2.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X582 XA8.XA12.MP0.G XA8.XA11.MN1.G XA8.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X583 AVSS XA6.XA4.MN0.G XA6.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X584 SARN XA0.XA11.MN1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X585 AVDD XA0.XA6.MP0.G XA0.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X586 VREF XA2.XA1.XA5.MN2.D XA2.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R74 XDAC1.XC0.XRES8.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X587 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X588 XA5.XA4.MN0.G XA5.XA1.XA5.MN2.G XA5.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X589 XA8.XA7.MP0.D XA8.XA7.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R75 D<8> XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X590 AVSS XA6.XA3.MN0.G D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X591 AVSS XA0.XA1.XA5.MN2.D D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X592 XA2.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X593 XA5.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X594 XA4.XA11.MN1.G XA3.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X595 AVSS XA20.XA2a.MN0.D XA1.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X596 XA1.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA1.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X597 XA4.XA11.MN1.G XA3.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X598 XA2.XA4.MN0.D XA2.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X599 XA0.XA1.XA4.MN1.D XA0.XA1.XA2.MP0.D XA0.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X600 XA4.XA8.MP0.D XA4.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X601 XA8.XA11.MP0.D XA8.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R76 m3_n2104_132# XB1.XA4.MP0.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X602 XA4.XA6.MP0.G XA4.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X603 XA0.XA6.MP2.G D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X604 XA0.XA1.XA1.MN0.D EN XA0.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X605 XA6.XA9.MN1.G CK_SAMPLE XA6.XA6.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X606 SARP XA0.XA11.MN1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X607 D<8> XA0.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X608 AVSS XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X609 VREF XA1.XA4.MN0.D XA1.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X610 AVSS XA1.XA4.MN0.D XA1.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X611 VREF XA7.XA1.XA5.MN2.D XA7.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R77 XDAC1.XC128b<2>.XRES1A.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X612 XA0.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X613 XA2.XA10.MP0.D XA2.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X614 AVSS XA1.XA3.MN0.G D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R78 m3_16472_308# XB2.XA3.MN1.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X615 XA7.XA1.XA4.MN1.D XA7.XA1.XA2.MP0.D XA7.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X616 VREF XA1.XA3.MN0.G D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X617 AVSS XA20.XA2a.MN0.D XA5.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X618 XA7.XA1.XA4.MP1.D EN XA7.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X619 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X620 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X621 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X622 AVSS XA6.XA11.MN1.G XA6.XA12.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X623 D<1> XA7.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X624 XA2.XA6.MP2.D D<6> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X625 D<1> XA7.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X626 XA7.XA1.XA1.MN0.D XA7.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X627 AVDD EN XA7.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X628 XA3.XA9.MN0.D XA3.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X629 XA6.XA4.MN0.G EN XA6.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X630 XA3.XA10.MP0.G XA3.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X631 XA6.XA7.MP0.D XA7.XA1.XA5.MN2.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X632 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R79 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X633 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X634 XA6.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA7.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X635 AVDD XA2.XA9.MN1.G XA2.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X636 XA1.XA6.MP0.G XA1.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X637 AVSS XA5.XA4.MN0.D XA5.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X638 XA7.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X639 XA1.XA6.MP0.G XA1.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X640 XA7.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X641 XA0.XA8.MP0.D XA0.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X642 XA6.XA12.MP0.G XA6.XA10.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X643 AVDD XA2.XA6.MP0.G XA2.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X644 XA8.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X645 AVSS XA5.XA3.MN0.G D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X646 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X647 XA0.XA6.MP0.G XA0.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X648 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X649 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X650 XB2.XA4.MP0.D XB2.XA0.MP0.D XB2.M1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X651 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X652 XA2.XA4.MN0.G XA2.XA1.XA5.MN2.G XA2.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X653 XA4.XA6.MP0.D XA4.XA6.MP0.G XA4.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X654 XA2.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X655 XB2.XA4.MN0.D XB2.XA0.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X656 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X657 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X658 AVSS XA8.XA4.MN0.D XA8.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X659 XA6.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA6.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X660 XA7.XA8.MP0.D XA7.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X661 XA5.XA6.MP0.G XA5.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X662 XB1.XA1.MN0.D XB1.XA1.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X663 XA7.XA8.MP0.D XA7.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R80 XDAC1.XC64a<0>.XRES4.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R81 XDAC1.XC0.XRES1A.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X664 SAR_IN XB2.XA0.MP0.D XB2.XA3.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X665 XA7.XA6.MP0.G XA7.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X666 AVSS XA8.XA4.MN0.G XA8.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X667 XA2.XA11.MN1.G XA1.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X668 XA7.XA6.MP0.G XA7.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X669 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X670 XA2.XA11.MN1.G XA1.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X671 VREF XA4.XA4.MN0.D XA4.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R82 XDAC1.X16ab.XRES16.B XA2.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X672 AVSS XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X673 SAR_IN XB2.XA3.MN0.S XB2.XA3.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X674 VREF XA6.XA4.MN0.D XA6.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X675 VREF XA4.XA4.MN0.G XA4.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R83 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X676 XB1.M1.G XB1.XA1.MP0.D XB1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X677 AVSS XA20.XA2a.MN0.D XA2.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X678 XA8.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X679 VREF XA6.XA3.MN0.G D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X680 VREF XA4.XA1.XA5.MN2.D XA4.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R84 XDAC1.XC64b<1>.XRES16.B D<7> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R85 XB1.XA3.MN1.D m3_7544_2420# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X681 XA8.XA4.MN0.D XA8.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X682 VREF XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R86 XA3.XA3.MN0.G XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X683 XA4.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X684 XA6.XA11.MN1.G XA5.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X685 XA5.XA1.XA4.MP1.D EN XA5.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X686 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X687 XA20.XA2.MN1.D SARP XA20.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X688 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X689 AVSS XA2.XA4.MN0.D XA2.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X690 XA4.XA4.MN0.D XA4.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X691 XA20.XA3a.MN0.G XA20.XA9.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R87 D<8> XDAC2.XC128a<1>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X692 SARN XB2.M1.G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X693 D<3> XA5.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X694 AVSS XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R88 XDAC1.XC64a<0>.XRES16.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X695 AVDD EN XA5.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X696 XA1.XA9.MN0.D XA1.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X697 XA6.XA6.MP0.G XA6.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X698 AVDD XA20.XA3a.MN0.G XA20.XA3a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X699 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X700 XA1.XA10.MP0.G XA1.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X701 AVSS XA2.XA3.MN0.G D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X702 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X703 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X704 XA8.XA10.MP0.D XA8.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X705 AVSS XA20.XA3.MN6.D XA20.XA2a.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X706 AVDD XA20.XA3.MN6.D XA20.XA2a.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X707 XA0.XA1.XA5.MN2.D EN XA0.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R89 XDAC1.XC0.XRES1B.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X708 XA5.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X709 XA8.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X710 XA0.XA4.MN0.D XA0.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R90 m3_16472_2420# XB2.XA3.MN1.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X711 XA20.XA3.MN0.D SARP XA20.XA2.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R91 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X712 XA0.XA1.XA2.MP0.D XA0.XA7.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X713 AVDD AVDD XA20.XA2.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X714 XA4.XA10.MP0.D XA4.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X715 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X716 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X717 XA0.XA6.MP2.G D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X718 XA20.XA1.MN0.D SARP XA20.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X719 XA2.XA6.MP0.G XA2.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X720 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X721 XA4.XA6.MP2.D D<4> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X722 XA8.XA10.MP0.G XA8.XA9.MN1.G XA8.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X723 XA5.XA9.MN0.D XA5.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X724 XA20.XA3.MN0.D XA20.XA9.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X725 AVDD XA20.XA9.MP0.D XA20.XA3.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X726 XA0.XA1.XA5.MP1.D EN XA0.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R92 XA4.XA6.MP0.G XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X727 XB1.XA4.MP0.D XB1.XA0.MP0.D XB1.M1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X728 AVSS CK_SAMPLE XA8.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X729 VREF XA8.XA1.XA5.MN2.D XA8.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X730 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R93 XDAC1.XC1.XRES16.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X731 XA7.XA11.MN1.G XA6.XA12.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X732 AVDD XA4.XA9.MN1.G XA4.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X733 XA20.XA2a.MN0.D XA20.XA3.MN6.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X734 AVDD XA0.XA1.XA1.MN0.S XA0.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R94 m3_n2104_3300# XB1.XA4.MP0.D sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X735 XA5.XA8.MP0.D XA5.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X736 XA3.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X737 XA8.XA1.XA4.MP1.D EN XA8.XA1.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X738 XA3.XA6.MP0.D XA3.XA6.MP0.G XA3.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X739 VREF XA0.XA4.MN0.G XA0.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X740 AVDD XA4.XA6.MP0.G XA4.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X741 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X742 XA5.XA6.MP0.G XA5.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X743 D<0> XA8.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X744 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R95 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X745 AVDD EN XA8.XA1.XA1.MN0.S AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X746 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X747 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X748 VREF D<8> XA0.XA6.MP2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X749 XA4.XA4.MN0.G XA4.XA1.XA5.MN2.G XA4.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X750 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X751 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X752 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X753 XB1.XA0.MP0.D CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X754 SAR_IP XB1.XA0.MP0.D XB1.XA3.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X755 XA4.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X756 XA3.XA11.MN1.G XA2.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X757 XA8.XA1.XA4.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X758 AVSS XA3.XA4.MN0.D XA3.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X759 VREF XA3.XA4.MN0.D XA3.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X760 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X761 XA0.XA9.MN1.G XA0.XA6.MP2.G XA0.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X762 AVSS XA3.XA4.MN0.G XA3.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R96 XDAC1.XC32a<0>.XRES2.B D<2> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X763 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X764 VREF XA3.XA4.MN0.G XA3.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R97 XDAC2.XC32a<0>.XRES1A.A AVSS sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X765 XA20.XA10.MN0.D XA20.XA11.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X766 XA20.XA10.MN1.D XA20.XA11.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X767 XA6.XA10.MP0.G XA6.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X768 XA2.XA1.XA5.MN2.D EN XA2.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X769 AVSS XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X770 VREF XA3.XA1.XA5.MN2.D XA3.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X771 AVSS XA6.XA1.XA5.MN2.D XA6.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R98 XA3.XA3.MN0.G XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X772 XA20.XA4.MN0.D SARN XA20.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X773 XA2.XA4.MN0.D XA2.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X774 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R99 XDAC1.XC128a<1>.XRES2.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X775 XA2.XA1.XA2.MP0.D XA3.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R100 D<8> XDAC2.XC128a<1>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R101 XA0.XA6.MP0.G XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X776 XA3.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X777 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X778 XA6.XA1.XA4.MN1.D XA6.XA1.XA2.MP0.D XA6.XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X779 XA3.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X780 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X781 XA0.XA12.MP0.G XA0.XA11.MN1.G XA0.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X782 D<6> XA2.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X783 AVSS XA20.XA2a.MN0.D XA4.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X784 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X785 DONE XA8.XA7.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X786 XA3.XA4.MN0.D XA3.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X787 XA3.XA4.MN0.D XA3.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X788 D<2> XA6.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R102 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X789 XA20.XA9.MP0.D XA20.XA10.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X790 XA6.XA1.XA1.MN0.D XA6.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X791 XA20.XA9.MP0.D XA20.XA10.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X792 XA0.XA7.MP0.D XA0.XA7.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X793 XA8.XA6.MP0.G XA8.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X794 XA2.XA1.XA5.MP1.D EN XA2.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X795 XA2.XA9.MN0.D XA2.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X796 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X797 SARP XB1.M1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X798 XA0.XA4.MN0.G EN XA0.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X799 AVDD XA2.XA1.XA1.MN0.S XA2.XA1.XA1.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R103 XDAC1.XC64a<0>.XRES2.B XA1.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X800 AVSS XA4.XA4.MN0.D XA4.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X801 XA0.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X802 XA6.XA1.XA4.MN0.D XA20.XA2a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X803 XA0.XA11.MP0.D XA0.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X804 VREF XA2.XA4.MN0.G XA2.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X805 XA3.XA10.MP0.D XA3.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R104 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X806 XA3.XA10.MP0.D XA3.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X807 AVSS XA4.XA3.MN0.G D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X808 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X809 VREF XA2.XA3.MN0.G D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R105 XDAC1.X16ab.XRES8.B XA3.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X810 XA3.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X811 XA3.XA6.MP2.D D<5> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R106 XA7.XA6.MP0.G XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X812 XA1.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X813 XA7.XA4.MN0.G XA7.XA1.XA5.MN2.G XA7.XA1.XA4.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X814 XA1.XA6.MP0.D XA1.XA6.MP0.G XA1.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X815 XA7.XA4.MN0.G EN XA7.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X816 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X817 XA7.XA1.XA1.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X818 XA2.XA9.MN1.G D<6> XA2.XA6.MP2.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X819 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X820 XA7.XA1.XA1.MP1.D XA20.XA3a.MN0.D XA8.XA1.XA5.MN2.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X821 XA3.XA10.MP0.G XA3.XA9.MN1.G XA3.XA9.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X822 AVDD XA3.XA9.MN1.G XA3.XA10.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X823 XA6.XA8.MP0.D XA6.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X824 XA4.XA6.MP0.G XA4.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R107 D<8> XDAC2.XC128a<1>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X825 AVSS XA20.XA2a.MN0.D XA0.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X826 AVSS CK_SAMPLE XA3.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X827 XA6.XA6.MP0.G XA6.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X828 AVDD XA3.XA6.MP0.G XA3.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X829 AVSS XA1.XA4.MN0.D XA1.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X830 VREF XA1.XA4.MN0.D XA1.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X831 XA5.XA6.MN0.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X832 AVSS XA1.XA4.MN0.G XA1.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R108 XDAC1.XC128b<2>.XRES8.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X833 XA2.XA12.MP0.G XA2.XA11.MN1.G XA2.XA11.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X834 VREF XA1.XA4.MN0.G XA1.XA4.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R109 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X835 AVSS XA0.XA4.MN0.D XA0.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X836 XA2.XA7.MP0.D XA3.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X837 AVSS XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X838 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X839 AVSS XA20.XA2a.MN0.D XA7.XA1.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X840 AVSS D<8> XA0.XA6.MP2.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X841 VREF XA1.XA1.XA5.MN2.D XA1.XA3.MN0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X842 XA7.XA1.XA1.MP2.D XA20.XA2a.MN0.D XA7.XA1.XA1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X843 XA1.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R110 XB2.XA4.MP0.D m3_26048_1188# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X844 XA1.XA1.XA5.MP0.D EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X845 XA5.XA11.MN1.G XA4.XA12.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X846 XA2.XA11.MP0.D XA2.XA10.MP0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X847 AVSS XA5.XA4.MN0.D XA5.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X848 XA1.XA4.MN0.D XA1.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X849 XA8.XA1.XA5.MN2.D XA8.XA1.XA5.MN2.G XA8.XA1.XA5.MN1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R111 XDAC1.XC128a<1>.XRES4.B XA0.XA6.MP2.G sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
R112 XB2.XA4.MP0.D m3_26048_4356# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X850 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X851 XA1.XA4.MN0.D XA1.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X852 AVSS XA7.XA4.MN0.D XA7.XA6.MP0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X853 XA8.XA4.MN0.D XA8.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X854 VREF XA7.XA4.MN0.D XA7.XA6.MP0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X855 AVSS XA5.XA4.MN0.G XA5.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X856 XA8.XA1.XA2.MP0.D XA8.XA7.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X857 XA0.XA6.MP0.G XA0.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R113 XDAC1.XC1.XRES8.B XA0.XA4.MN0.D sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X858 XA4.XA1.XA5.MN2.D EN XA4.XA1.XA5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X859 AVSS XA7.XA3.MN0.G D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X860 D<0> XA8.XA3.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X861 VREF XA7.XA3.MN0.G D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X862 AVSS XA5.XA1.XA5.MN2.D XA5.XA3.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X863 XA4.XA4.MN0.D XA4.XA4.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R114 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X864 XA4.XA1.XA2.MP0.D XA5.XA1.XA5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X865 SARP XB1.M1.G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X866 XA5.XA1.XA5.MN0.D XA20.XA3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X867 XA8.XA1.XA5.MN1.D XA8.XA1.XA2.MP0.D XA8.XA1.XA5.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X868 XA1.XA10.MP0.D XA1.XA10.MP0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X869 XA1.XA10.MP0.D XA1.XA10.MP0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X870 XA6.XA6.MP0.D XA6.XA6.MP0.G XA6.XA9.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X871 D<4> XA4.XA3.MN0.G VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X872 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X873 XA5.XA4.MN0.D XA5.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X874 XA0.XA11.MN1.G XB1.XA2.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X875 XA8.XA7.MP0.G XA8.XA1.XA1.MN0.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X876 XA1.XA6.MN2.D CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X877 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X878 XA1.XA6.MP2.D D<7> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X879 XA4.XA1.XA5.MP1.D EN XA4.XA1.XA5.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X880 XA4.XA9.MN0.D XA4.XA7.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X881 XA7.XA6.MP0.G XA7.XA4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X882 AVSS XA8.XA4.MN0.G XA8.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X883 XA7.XA6.MP0.G XA7.XA4.MN0.D VREF AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R115 XDAC1.XC32a<0>.XRES4.B D<3> sky130_fd_pr__res_generic_l1 w=0.38 l=0.3
X884 XB1.XA3.MN1.D XB1.XA0.MP0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X885 XA5.XA4.MN0.G EN XA5.XA1.XA4.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 a_17408_50436# a_18560_50436# 0.00133f
C1 D<3> a_13520_50084# 5.7e-19
C2 AVDD a_16040_45156# 0.356f
C3 D<7> a_2288_49732# 0.0109f
C4 XA7.XA1.XA5.MN2.G XA7.XA4.MN0.D 6.95e-19
C5 XA8.XA1.XA5.MN2.G XA6.XA4.MN0.D 6.95e-19
C6 XA6.XA1.XA4.MP1.D a_16040_42692# 0.049f
C7 XA1.XA1.XA4.MN1.D XA1.XA1.XA4.MN0.D 0.0488f
C8 VREF a_9848_48676# 1.3e-19
C9 AVDD a_23600_42692# 0.0232f
C10 XA2.XA6.MP0.G a_4808_47620# 4.4e-19
C11 XA6.XA6.MP0.G a_16040_47972# 8.92e-19
C12 D<3> XA2.XA3.MN0.G 0.0338f
C13 AVDD a_22448_54308# 0.364f
C14 XA5.XA1.XA1.MN0.S XA6.XA1.XA1.MN0.S 0.00217f
C15 XA1.XA1.XA1.MN0.S a_2288_41284# 0.0948f
C16 a_14888_41636# a_14888_41284# 0.0109f
C17 XA0.XA6.MP0.G a_920_44100# 5.5e-19
C18 XA4.XA1.XA5.MN2.G a_9848_43396# 0.00504f
C19 a_18560_47620# a_19928_47620# 8.89e-19
C20 XA7.XA4.MN0.G a_17408_46916# 0.0662f
C21 XA4.XA6.MP0.G a_11000_44452# 5.5e-19
C22 VREF XA0.XA1.XA5.MN2.D 0.341f
C23 AVDD a_19928_39876# 0.00148f
C24 a_14888_53252# XA6.XA10.MP0.D 0.0692f
C25 a_4808_53252# a_4808_52900# 0.0109f
C26 AVDD a_14888_51844# 0.00166f
C27 XA7.XA11.MN1.G a_18560_52548# 0.00103f
C28 a_13520_40228# a_13520_39876# 0.0109f
C29 XA2.XA6.MP0.G a_4808_41988# 7.76e-20
C30 SARN a_14960_3854# 2.37e-19
C31 XA20.XA2a.MN0.D XA4.XA1.XA5.MN2.D 8.92e-20
C32 a_13520_45860# a_14888_45860# 8.89e-19
C33 XA6.XA6.MP0.G a_14888_42340# 7.76e-20
C34 XA4.XA4.MN0.G a_11000_43748# 6.3e-19
C35 XA1.XA3.MN0.G a_2288_44804# 0.00498f
C36 XA8.XA3.MN0.G a_19928_45156# 0.0805f
C37 XA20.XA3a.MN0.D XA1.XA1.XA5.MP1.D 2.15e-19
C38 XA4.XA1.XA5.MN2.G a_8480_40932# 0.00838f
C39 XA20.XA3.MN0.D a_23600_42692# 0.00454f
C40 XA3.XA9.MN1.G a_9848_51492# 2.84e-19
C41 XA1.XA7.MP0.D a_2288_51844# 0.133f
C42 AVDD XA8.XA4.MN0.D 2.57f
C43 CK_SAMPLE a_22448_50084# 5.94e-19
C44 XA7.XA4.MN0.G XA7.XA1.XA1.MN0.S 5.22e-20
C45 XA0.XA6.MP2.G li_9184_29616# 3.5e-20
C46 SARN XDAC2.XC32a<0>.XRES2.B 6.99f
C47 a_7328_44100# a_8480_44100# 0.00133f
C48 a_16040_44452# EN 0.00173f
C49 XA20.XA3a.MN0.D a_14888_41636# 0.00547f
C50 a_8480_45156# XA3.XA1.XA2.MP0.D 1.56e-20
C51 XA20.XA2a.MN0.D a_920_42692# 0.00457f
C52 XA7.XA9.MN1.G a_18560_49380# 4.23e-20
C53 AVDD a_13520_46212# 0.00125f
C54 D<7> a_2288_50436# 0.0863f
C55 D<3> a_12368_50788# 0.161f
C56 a_2288_51140# XA1.XA6.MP0.G 6.76e-20
C57 XDAC2.XC128a<1>.XRES8.B li_14804_17952# 9.91e-20
C58 XDAC1.XC128a<1>.XRES8.B XDAC1.XC128a<1>.XRES2.B 0.44f
C59 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES16.B 0.0483f
C60 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES1A.B 0.00438f
C61 XA8.XA1.XA2.MP0.D XA8.XA1.XA4.MN1.D 0.056f
C62 a_7328_43044# a_8480_43044# 0.00133f
C63 XA0.XA6.MP0.G li_14804_8736# 0.00506f
C64 EN a_2288_41988# 0.0723f
C65 D<7> a_3440_47620# 5.21e-19
C66 XA6.XA1.XA5.MN2.G a_12368_47268# 0.00363f
C67 AVDD a_7328_43396# 0.361f
C68 a_5960_49732# XA2.XA4.MN0.D 0.0658f
C69 a_18560_41988# a_19928_41988# 8.89e-19
C70 XA8.XA7.MP0.G a_22448_44100# 0.0012f
C71 AVDD a_5960_40932# 0.358f
C72 XA2.XA1.XA5.MN2.G XA2.XA1.XA5.MN1.D 0.0102f
C73 D<2> SARP 0.0407f
C74 XA7.XA1.XA5.MN2.G EN 0.946f
C75 XA4.XA6.MP0.G a_11000_45508# 5.5e-19
C76 VREF a_12368_46564# 0.0175f
C77 XA3.XA4.MN0.D a_8480_46564# 0.001f
C78 XA5.XA11.MN1.G a_9848_53252# 2.82e-19
C79 DONE XA20.XA4.MN0.D 0.00191f
C80 a_16040_53604# a_17408_53604# 8.89e-19
C81 AVDD a_11000_52548# 0.405f
C82 a_5960_40580# a_7328_40580# 8.89e-19
C83 XA3.XA6.MP0.G XA3.XA1.XA4.MN1.D 7.41e-19
C84 XA6.XA1.XA5.MN2.G a_12368_41636# 0.0736f
C85 XA5.XA1.XA5.MN2.G a_13520_41636# 0.0039f
C86 D<7> a_3440_41988# 6.49e-19
C87 XA7.XA3.MN0.G a_18560_46212# 0.157f
C88 XA0.XA4.MN0.G a_920_44452# 5.54e-19
C89 XA7.XA4.MN0.G a_18560_44804# 0.00858f
C90 XA7.XA6.MP0.G a_18560_43044# 7.76e-20
C91 XA0.XA11.MN1.G XB2.XA0.MP0.D 0.0801f
C92 D<3> a_13520_42340# 6.49e-19
C93 AVDD XA3.XA6.MP0.G 5.93f
C94 XA0.XA10.MP0.G a_920_51844# 0.00224f
C95 XA5.XA10.MP0.G XA5.XA7.MP0.D 0.0601f
C96 a_n232_52548# XA0.XA7.MP0.D 5.16e-20
C97 CK_SAMPLE a_21080_50788# 0.00554f
C98 a_12368_52548# a_12368_52196# 0.0109f
C99 XA0.XA9.MN1.G a_n232_52196# 0.0862f
C100 SAR_IN a_13808_334# 1.73e-19
C101 XA20.XA3a.MN0.D XA0.XA1.XA4.MN0.D 1.1e-19
C102 XA20.XA2a.MN0.D XA5.XA1.XA2.MP0.D 0.227f
C103 XA3.XA6.MP0.G a_7328_40228# 2.44e-19
C104 XA3.XA4.MN0.G a_8480_42340# 7.97e-19
C105 XA4.XA1.XA5.MN2.D a_11000_44100# 0.126f
C106 a_16040_45508# EN 1.42e-19
C107 XA7.XA6.MP0.G a_17408_40580# 5.5e-19
C108 SARN XA7.XA6.MP0.G 0.0461f
C109 XA2.XA9.MN1.G a_5960_50084# 0.00281f
C110 a_n232_51140# XA0.XA6.MN2.D 0.00176f
C111 a_920_51140# XA0.XA6.MP2.G 0.0672f
C112 a_12368_51140# a_13520_51140# 0.00133f
C113 XA3.XA1.XA5.MN2.G XA2.XA6.MP2.D 0.00313f
C114 AVDD a_12368_47268# 0.356f
C115 a_21080_52900# VREF 0.00386f
C116 XB1.XA4.MP0.D m3_n1960_4356# 0.0137f
C117 EN XA4.XA1.XA4.MN1.D 3.17e-19
C118 XA20.XA2a.MN0.D XA2.XA1.XA1.MP1.D 0.00946f
C119 XA1.XA6.MN0.D a_3440_49732# 0.00176f
C120 AVDD XA0.XA1.XA5.MN1.D 0.00889f
C121 D<3> a_12368_49028# 0.00884f
C122 D<7> a_2288_48676# 0.00918f
C123 XA5.XA1.XA5.MN2.G a_12368_48324# 7.1e-20
C124 XA6.XA1.XA5.MN2.G a_11000_48324# 7.1e-20
C125 D<8> XDAC2.X16ab.XRES2.B 4.06e-21
C126 a_11000_43044# XA4.XA1.XA1.MN0.S 4.06e-20
C127 D<1> a_19928_45860# 1.06e-19
C128 XA6.XA1.XA5.MN2.G a_14888_45156# 1e-19
C129 a_17408_48676# a_18560_48676# 0.00133f
C130 XA6.XA6.MP0.G XA2.XA3.MN0.G 0.21f
C131 XA20.XA10.MN1.D a_23600_42692# 0.00386f
C132 AVDD a_12368_41636# 0.404f
C133 VREF a_9848_47620# 7.12e-19
C134 XA2.XA6.MP0.G a_5960_46564# 5.5e-19
C135 XA5.XA6.MP0.G XA5.XA3.MN0.G 0.05f
C136 XA20.XA11.MN0.D a_23600_53604# 0.0949f
C137 DONE a_22448_53604# 0.006f
C138 AVDD XA7.XA11.MP0.D 0.176f
C139 a_22448_54308# XA20.XA10.MN1.D 1.28e-19
C140 a_8480_53956# XA3.XA12.MP0.G 0.0688f
C141 a_9848_53956# XA4.XA11.MN1.G 7.59e-19
C142 a_11000_41284# a_11000_40932# 0.0109f
C143 XA4.XA1.XA1.MN0.S a_9848_40580# 0.00155f
C144 XA0.XA4.MN0.D a_n232_44100# 9.25e-20
C145 XA2.XA6.MP0.G XA2.XA1.XA2.MP0.D 0.0106f
C146 XA0.XA4.MN0.G a_920_45508# 6.57e-19
C147 XA7.XA4.MN0.G a_17408_45860# 2.12e-19
C148 AVDD a_13808_1038# 0.00181f
C149 a_12368_46916# a_13520_46916# 0.00133f
C150 a_920_46916# D<8> 0.0658f
C151 XA8.XA1.XA5.MN2.G a_19928_42692# 0.0739f
C152 XA2.XA1.XA5.MN2.G XA1.XA1.XA4.MP0.D 0.00361f
C153 XA0.XA7.MP0.G XA1.XA1.XA4.MN0.D 0.00313f
C154 XA4.XA11.MN1.G XA3.XA8.MP0.D 2.37e-19
C155 a_11000_52900# a_11000_52548# 0.0109f
C156 a_23600_52900# XA20.XA4.MN0.D 0.00176f
C157 XA20.XA9.MP0.D a_23600_52548# 0.0765f
C158 XA8.XA11.MN1.G a_18560_51844# 1.13e-19
C159 AVDD XA1.XA6.MN2.D 3.77e-19
C160 CK_SAMPLE XA3.XA1.XA5.MN2.G 0.0595f
C161 a_14960_3150# a_14960_2798# 0.0109f
C162 a_13808_3854# XB2.XA1.MP0.D 1.01e-19
C163 XA5.XA4.MN0.G a_13520_43044# 0.0409f
C164 XA7.XA1.XA5.MN2.G a_17408_39876# 0.00278f
C165 D<6> a_5960_40228# 7.76e-20
C166 D<2> a_16040_40580# 4.07e-20
C167 SARN a_12368_334# 0.0348f
C168 XA20.XA3a.MN0.D a_8480_43396# 0.0723f
C169 XA6.XA1.XA5.MN2.D XA7.XA1.XA5.MN2.D 0.00869f
C170 XA1.XA1.XA5.MN2.D a_3440_45156# 0.153f
C171 a_14888_45508# a_14888_45156# 0.0109f
C172 XA5.XA8.MP0.D a_13520_51492# 0.00224f
C173 a_22448_51844# a_22448_51492# 0.0109f
C174 XA7.XA9.MN1.G D<1> 0.0378f
C175 XA5.XA7.MP0.D a_13520_51140# 0.00388f
C176 AVDD a_11000_48324# 0.359f
C177 XA2.XA9.MN1.G a_4808_50788# 0.015f
C178 a_7328_53604# VREF 0.00396f
C179 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES16.B 0.0483f
C180 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES1A.B 0.00438f
C181 XDAC2.XC64b<1>.XRES8.B XDAC2.XC64b<1>.XRES2.B 0.44f
C182 XA20.XA3a.MN0.D a_7328_40932# 0.0674f
C183 XA20.XA2a.MN0.D a_14888_41988# 0.0844f
C184 XA20.XA2.MN1.D a_23600_43044# 0.00245f
C185 a_2288_43748# a_3440_43748# 0.00133f
C186 XA0.XA6.MP2.G XDAC1.XC128a<1>.XRES1B.B 0.00406f
C187 EN XA1.XA1.XA5.MP0.D 0.0446f
C188 XA0.XA1.XA5.MP1.D XA0.XA1.XA5.MP0.D 0.0488f
C189 D<3> a_12368_50084# 0.0155f
C190 AVDD a_14888_45156# 0.00125f
C191 a_3440_50436# XA1.XA6.MN0.D 0.00176f
C192 XA7.XA1.XA5.MN2.G XA6.XA4.MN0.D 0.0939f
C193 XA2.XA1.XA5.MN2.G a_2288_49380# 0.00363f
C194 XDAC2.XC32a<0>.XRES8.B XDAC2.XC64a<0>.XRES8.B 6.7e-19
C195 li_14804_13248# li_14804_12636# 0.00271f
C196 a_3440_42692# a_4808_42692# 8.89e-19
C197 XA6.XA1.XA4.MN1.D a_16040_42692# 2.16e-19
C198 XA6.XA1.XA4.MP1.D a_14888_42692# 2.16e-19
C199 EN a_17408_41284# 0.00564f
C200 XA0.XA4.MN0.D li_9184_8736# 0.00506f
C201 VREF a_8480_48676# 1.3e-19
C202 XA2.XA4.MN0.D a_5960_48676# 0.154f
C203 AVDD a_22448_42692# 0.471f
C204 XA6.XA6.MP0.G a_14888_47972# 6.28e-19
C205 D<3> XA1.XA3.MN0.G 0.0259f
C206 a_11000_49380# a_11000_49028# 0.0109f
C207 XA6.XA1.XA5.MN2.G a_12368_46212# 0.00363f
C208 D<4> XA4.XA3.MN0.G 0.572f
C209 D<1> a_18560_46916# 0.00249f
C210 AVDD a_21080_54308# 0.447f
C211 a_2288_54308# a_3440_54308# 0.00133f
C212 SARP li_9184_24300# 0.00103f
C213 XA5.XA1.XA1.MN0.S XA5.XA1.XA1.MP2.D 0.0708f
C214 XA4.XA1.XA5.MN2.G a_8480_43396# 2.66e-19
C215 XA3.XA1.XA5.MN2.G a_9848_43396# 7.1e-20
C216 D<7> XA1.XA1.XA5.MN0.D 0.00188f
C217 a_5960_47620# a_5960_47268# 0.0109f
C218 XA0.XA4.MN0.G D<8> 0.622f
C219 XA4.XA6.MP0.G a_9848_44452# 7.76e-20
C220 XA0.XA4.MN0.D XA0.XA1.XA5.MN2.D 0.0265f
C221 XA7.XA6.MP0.G SARP 0.029f
C222 AVDD a_18560_39876# 0.00131f
C223 XA0.XA6.MP0.G a_n232_44100# 7.76e-20
C224 XA2.XA11.MN1.G XA2.XA9.MN1.G 0.00804f
C225 a_22448_53252# a_23600_53252# 0.00133f
C226 AVDD a_13520_51844# 0.00166f
C227 XA7.XA11.MN1.G a_17408_52548# 0.00135f
C228 a_n232_39876# a_920_39876# 0.00133f
C229 SARN a_13808_3854# 0.00146f
C230 XA20.XA2a.MN0.D XA3.XA1.XA5.MN2.D 8.92e-20
C231 a_920_45860# a_920_45508# 0.0109f
C232 XA4.XA4.MN0.G a_9848_43748# 0.0157f
C233 XA20.XA3a.MN0.D XA0.XA1.XA5.MP1.D 2.15e-19
C234 XA3.XA1.XA5.MN2.G a_8480_40932# 0.00631f
C235 XA4.XA1.XA5.MN2.G a_7328_40932# 0.0245f
C236 XA20.XA3.MN0.D a_22448_42692# 0.0215f
C237 a_13520_52196# a_13520_51844# 0.0109f
C238 XA3.XA9.MN1.G a_8480_51492# 0.0118f
C239 a_22448_54660# VREF 0.00135f
C240 a_11000_52548# XA5.XA1.XA5.MN2.G 1.75e-19
C241 XA7.XA9.MN1.G XA7.XA8.MP0.D 0.0132f
C242 XA5.XA7.MP0.D XA6.XA7.MP0.D 0.00435f
C243 AVDD XA7.XA4.MN0.D 2.51f
C244 CK_SAMPLE a_21080_50084# 9.85e-19
C245 a_19928_44452# a_19928_44100# 0.0109f
C246 a_14888_44452# EN 0.00154f
C247 XA20.XA3a.MN0.D a_13520_41636# 0.00547f
C248 XA6.XA1.XA5.MN2.D XA6.XA1.XA2.MP0.D 4.72e-19
C249 XA20.XA2a.MN0.D a_n232_42692# 0.00563f
C250 a_22448_52196# VREF 0.00104f
C251 XA20.XA9.MP0.D a_23600_48324# 0.0714f
C252 AVDD a_12368_46212# 0.356f
C253 XA7.XA9.MN1.G a_17408_49380# 2.54e-19
C254 XA4.XA1.XA2.MP0.D a_11000_42692# 7.68e-20
C255 XA0.XA1.XA2.MP0.D XA0.XA1.XA4.MP0.D 4.34e-19
C256 a_19928_43396# a_19928_43044# 0.0109f
C257 EN a_920_41988# 0.0739f
C258 XA1.XA6.MP0.G li_14804_9156# 0.00504f
C259 D<6> XA20.XA3a.MN0.D 0.0701f
C260 D<7> a_2288_47620# 0.0147f
C261 XA5.XA1.XA5.MN2.G a_12368_47268# 7.1e-20
C262 XA6.XA1.XA5.MN2.G a_11000_47268# 7.1e-20
C263 AVDD a_5960_43396# 0.361f
C264 D<3> a_13520_47972# 5.43e-19
C265 XA20.XA3.MN1.D a_23600_49380# 0.0605f
C266 a_16040_49732# a_17408_49732# 8.89e-19
C267 a_4808_49732# XA2.XA4.MN0.D 0.0675f
C268 a_7328_49732# VREF 0.029f
C269 a_5960_41988# a_5960_41636# 0.0109f
C270 XA6.XA1.XA5.MN2.G EN 0.897f
C271 D<5> a_8480_44452# 5.26e-19
C272 XA8.XA7.MP0.G a_21080_44100# 0.00556f
C273 AVDD a_4808_40932# 0.00125f
C274 XA2.XA1.XA5.MN2.G XA1.XA1.XA5.MN1.D 6.68e-19
C275 XA0.XA6.MP0.G XA0.XA1.XA5.MN2.D 0.0268f
C276 a_n232_47972# a_920_47972# 0.00133f
C277 XA3.XA4.MN0.G a_8480_47972# 0.153f
C278 a_18560_48324# a_18560_47972# 0.0109f
C279 XA4.XA6.MP0.G a_9848_45508# 7.76e-20
C280 VREF a_11000_46564# 0.0175f
C281 XA3.XA4.MN0.D a_7328_46564# 2.2e-19
C282 XA4.XA11.MN1.G a_11000_53252# 0.0674f
C283 DONE XA8.XA10.MP0.G 0.0577f
C284 XA8.XA12.MP0.G XA8.XA11.MP0.D 0.0612f
C285 AVDD a_9848_52548# 0.00166f
C286 a_18560_40932# a_18560_40580# 0.0109f
C287 XA7.XA3.MN0.G a_17408_46212# 0.155f
C288 D<8> a_920_45860# 0.155f
C289 XA7.XA4.MN0.G a_17408_44804# 5.54e-19
C290 XA0.XA4.MN0.G a_n232_44452# 0.00907f
C291 XA3.XA6.MP0.G XA3.XA1.XA4.MP1.D 0.00121f
C292 XA5.XA1.XA5.MN2.G a_12368_41636# 4.13e-19
C293 D<7> a_2288_41988# 7.77e-20
C294 XA7.XA6.MP0.G a_17408_43044# 5.5e-19
C295 XA2.XA4.MN0.D XA2.XA1.XA5.MP0.D 9.69e-19
C296 VREF XA3.XA1.XA5.MP0.D 0.00202f
C297 XA0.XA11.MN1.G XB1.XA0.MP0.D 0.0801f
C298 a_19928_46564# a_21080_46564# 0.00133f
C299 a_7328_46564# a_7328_46212# 0.0109f
C300 D<3> a_12368_42340# 7.77e-20
C301 AVDD XA2.XA6.MP0.D 0.144f
C302 XA0.XA10.MP0.G a_n232_51844# 5.59e-19
C303 CK_SAMPLE a_19928_50788# 0.164f
C304 XA4.XA9.MN1.G XA5.XA9.MN1.G 0.00217f
C305 XB2.M1.G a_14960_1038# 1.7e-19
C306 SAR_IN a_12368_334# 0.0566f
C307 XB1.M1.G a_11000_686# 0.161f
C308 a_8408_1742# a_8408_1390# 0.0109f
C309 a_13520_44804# a_14888_44804# 8.89e-19
C310 a_920_44804# a_920_44452# 0.0109f
C311 XA3.XA4.MN0.G a_7328_42340# 1.28e-19
C312 XA5.XA3.MN0.G a_13520_43396# 6.8e-20
C313 XA4.XA1.XA5.MN2.D a_9848_44100# 0.0877f
C314 a_14888_45508# EN 3.34e-19
C315 XA7.XA6.MP0.G a_16040_40580# 1.36e-19
C316 SARN XDAC2.X16ab.XRES2.B 6.99f
C317 XA2.XA9.MN1.G a_4808_50084# 0.00969f
C318 XA4.XA1.XA5.MN2.G D<6> 3.47e-19
C319 XA3.XA1.XA5.MN2.G XA2.XA6.MN2.D 6.33e-19
C320 AVDD a_11000_47268# 0.356f
C321 XB1.XA4.MP0.D m3_n2104_4356# 0.0273f
C322 XDAC1.X16ab.XRES1A.B XDAC1.XC128b<2>.XRES1B.B 0.617f
C323 EN XA3.XA1.XA4.MN1.D 3.17e-19
C324 XA20.XA2a.MN0.D XA2.XA1.XA1.MN0.D 0.0221f
C325 XA1.XA1.XA5.MN0.D a_3440_43396# 0.0474f
C326 a_17408_43748# a_17408_43396# 0.0109f
C327 XA5.XA6.MN0.D a_13520_50084# 0.0488f
C328 AVDD EN 40.3f
C329 a_7328_50436# VREF 0.0035f
C330 XA5.XA1.XA5.MN2.G a_11000_48324# 0.00455f
C331 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES2.B 0.0307f
C332 li_9184_8124# li_9184_7512# 0.00271f
C333 XDAC1.XC64a<0>.XRES1A.B XDAC1.XC1.XRES1A.B 0.00444f
C334 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES16.B 0.0381f
C335 XA3.XA3.MN0.G XDAC2.X16ab.XRES8.B 1.85e-19
C336 XA4.XA1.XA4.MP0.D a_11000_42340# 0.049f
C337 a_23600_42692# a_23600_42340# 0.0109f
C338 EN a_7328_40228# 0.0658f
C339 D<1> a_18560_45860# 0.0675f
C340 XA6.XA1.XA5.MN2.G a_13520_45156# 1.95e-19
C341 a_4808_48676# a_4808_48324# 0.0109f
C342 XA6.XA6.MP0.G XA1.XA3.MN0.G 0.0265f
C343 AVDD a_11000_41636# 0.404f
C344 XA2.XA4.MN0.D a_5960_47620# 0.00498f
C345 VREF a_8480_47620# 7.12e-19
C346 D<5> a_8480_45508# 0.0031f
C347 XA2.XA6.MP0.G a_4808_46564# 7.76e-20
C348 XA20.XA11.MN0.D a_22448_53604# 0.0674f
C349 DONE a_21080_53604# 0.00126f
C350 AVDD XA6.XA11.MP0.D 0.19f
C351 CK_SAMPLE XA8.XA11.MN1.G 0.0011f
C352 a_19928_53956# a_21080_53956# 0.00133f
C353 a_7328_53956# XA3.XA12.MP0.G 0.0674f
C354 a_8480_53956# XA4.XA11.MN1.G 0.0225f
C355 SARP XDAC1.XC32a<0>.XRES2.B 6.99f
C356 VREF a_22448_44452# 3.15e-19
C357 D<2> a_16040_43044# 7.76e-20
C358 XA6.XA6.MP0.G a_16040_43748# 5.5e-19
C359 XA0.XA4.MN0.G a_n232_45508# 0.0104f
C360 a_n232_46916# D<8> 0.0682f
C361 D<6> XA2.XA1.XA4.MP1.D 7.42e-19
C362 XA8.XA1.XA5.MN2.G a_18560_42692# 1.95e-19
C363 XA0.XA7.MP0.G XA1.XA1.XA4.MP0.D 6.33e-19
C364 XA3.XA10.MP0.G XA4.XA10.MP0.G 0.00217f
C365 AVDD XA1.XA6.MP2.D 0.172f
C366 CK_SAMPLE XA2.XA1.XA5.MN2.G 0.0595f
C367 a_9560_2798# a_11000_2798# 8e-19
C368 XA3.XA3.MN0.G XA3.XA1.XA5.MN1.D 0.00103f
C369 XA5.XA4.MN0.G a_12368_43044# 0.0222f
C370 XA7.XA1.XA5.MN2.G a_16040_39876# 0.00285f
C371 D<6> a_4808_40228# 6.49e-19
C372 XA4.XA6.MP0.G a_11000_41284# 4.24e-19
C373 XA2.XA4.MN0.D a_5960_41988# 9.14e-20
C374 D<2> a_14888_40580# 5.24e-19
C375 SARN a_11000_334# 2.76e-20
C376 XA20.XA3a.MN0.D a_7328_43396# 0.00213f
C377 XA1.XA1.XA5.MN2.D a_2288_45156# 0.155f
C378 AVDD a_9848_48324# 0.00131f
C379 XA5.XA8.MP0.D a_12368_51492# 0.00224f
C380 a_3440_51492# a_4808_51492# 8.89e-19
C381 a_12368_51844# XA6.XA1.XA5.MN2.G 8.87e-19
C382 XA5.XA7.MP0.D a_12368_51140# 0.00224f
C383 CK_SAMPLE a_19928_49028# 3.19e-19
C384 a_5960_53604# VREF 0.00351f
C385 a_7328_52196# D<5> 7.56e-20
C386 XA20.XA3a.MN0.D a_5960_40932# 0.0658f
C387 XA3.XA1.XA5.MN2.D a_7328_42692# 7.44e-20
C388 XA20.XA2a.MN0.D a_13520_41988# 0.0861f
C389 XA20.XA2.MN1.D a_22448_43044# 0.00245f
C390 XA5.XA1.XA5.MN1.D a_13520_43748# 0.0494f
C391 D<8> XA0.XA1.XA1.MN0.S 0.0101f
C392 EN XA1.XA1.XA2.MP0.D 0.03f
C393 a_16040_50436# a_17408_50436# 8.89e-19
C394 AVDD a_13520_45156# 0.00125f
C395 XA20.XA9.MP0.D a_23600_47268# 0.00334f
C396 a_2288_51140# VREF 0.00383f
C397 XA0.XA7.MP0.G a_2288_49380# 7.1e-20
C398 XA2.XA1.XA5.MN2.G a_920_49380# 7.1e-20
C399 EN a_16040_41284# 0.00564f
C400 XA1.XA1.XA4.MP1.D XA1.XA1.XA4.MP0.D 0.0488f
C401 XA6.XA1.XA4.MN1.D a_14888_42692# 0.0474f
C402 XA2.XA4.MN0.D a_4808_48676# 0.158f
C403 VREF a_7328_48676# 0.0191f
C404 XA3.XA6.MP0.G XA20.XA3a.MN0.D 0.0676f
C405 D<3> D<8> 0.0322f
C406 a_22448_49380# a_23600_49380# 0.00133f
C407 D<7> a_3440_46564# 0.0551f
C408 XA5.XA1.XA5.MN2.G a_12368_46212# 7.1e-20
C409 XA6.XA1.XA5.MN2.G a_11000_46212# 7.1e-20
C410 D<4> XA3.XA3.MN0.G 0.225f
C411 D<1> a_17408_46916# 0.0185f
C412 AVDD a_21080_42692# 0.359f
C413 AVDD a_19928_54308# 0.00166f
C414 XA0.XA1.XA1.MP2.D a_920_41284# 0.0465f
C415 a_13520_41636# a_13520_41284# 0.0109f
C416 XA4.XA1.XA5.MN2.G a_7328_43396# 0.00442f
C417 XA3.XA1.XA5.MN2.G a_8480_43396# 0.00518f
C418 D<7> XA1.XA1.XA5.MP0.D 7.43e-19
C419 a_17408_47620# a_18560_47620# 0.00133f
C420 XA6.XA4.MN0.G a_16040_46916# 0.0678f
C421 VREF a_22448_45508# 9.89e-19
C422 AVDD a_17408_39876# 0.438f
C423 XA5.XA11.MP0.D a_12368_52900# 0.00176f
C424 a_13520_53252# XA5.XA10.MP0.D 0.0676f
C425 a_3440_53252# a_3440_52900# 0.0109f
C426 AVDD a_12368_51844# 0.387f
C427 XA2.XA11.MN1.G XA1.XA9.MN0.D 1.71e-19
C428 XA7.XA11.MN1.G a_16040_52548# 9.29e-19
C429 a_12368_40228# a_12368_39876# 0.0109f
C430 XA20.XA2a.MN0.D XA2.XA1.XA5.MN2.D 8.92e-20
C431 a_12368_45860# a_13520_45860# 0.00133f
C432 D<8> a_920_44804# 0.00498f
C433 XA7.XA3.MN0.G a_18560_45156# 0.0805f
C434 XA20.XA3a.MN0.D XA0.XA1.XA5.MN1.D 2.15e-19
C435 XA3.XA1.XA5.MN2.G a_7328_40932# 0.0013f
C436 D<1> XA7.XA1.XA1.MN0.S 0.0159f
C437 XA3.XA9.MN1.G a_7328_51492# 6.57e-19
C438 XA20.XA12.MP0.G VREF 0.188f
C439 XA0.XA7.MP0.D a_920_51844# 0.133f
C440 AVDD XA6.XA4.MN0.D 2.51f
C441 CK_SAMPLE a_19928_50084# 0.162f
C442 XA0.XA6.MP2.G XDAC1.XC64b<1>.XRES1B.B 4.06e-21
C443 a_13520_44452# EN 0.00154f
C444 SARN li_14804_14472# 0.00103f
C445 a_5960_44100# a_7328_44100# 8.89e-19
C446 XA20.XA2a.MN0.D XA8.XA1.XA4.MP1.D 0.00728f
C447 XA4.XA6.MP2.D a_11000_50788# 0.049f
C448 a_21080_52196# VREF 0.00386f
C449 XA0.XA6.MP2.D a_920_50436# 0.00176f
C450 D<0> XA8.XA6.MP2.D 0.0399f
C451 XA4.XA1.XA5.MN2.G XA3.XA6.MP0.G 0.174f
C452 XA20.XA9.MP0.D a_22448_48324# 0.139f
C453 AVDD a_11000_46212# 0.356f
C454 XDAC1.XC128a<1>.XRES8.B li_9184_17952# 9.91e-20
C455 li_14804_18564# li_14804_17952# 0.00271f
C456 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES2.B 0.0307f
C457 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES16.B 0.0381f
C458 XDAC2.XC128b<2>.XRES1A.B XDAC2.XC128a<1>.XRES1A.B 0.00444f
C459 XA20.XA2a.MN0.D a_19928_40228# 2.1e-19
C460 XA0.XA1.XA2.MP0.D XA0.XA1.XA4.MN0.D 0.056f
C461 XA4.XA1.XA2.MP0.D a_9848_42692# 0.0962f
C462 a_5960_43044# a_7328_43044# 8.89e-19
C463 XA0.XA6.MP0.G XDAC2.XC1.XRES1B.B 0.00405f
C464 EN a_n232_41988# 0.00418f
C465 XA5.XA1.XA5.MN2.G a_11000_47268# 0.00363f
C466 AVDD a_4808_43396# 0.00125f
C467 XA20.XA10.MN1.D EN 0.00237f
C468 D<3> a_12368_47972# 0.0147f
C469 XA20.XA3.MN6.D a_23600_49380# 6.01e-19
C470 XA20.XA3.MN1.D a_22448_49380# 8.29e-20
C471 a_5960_49732# VREF 0.029f
C472 SARP a_11000_334# 0.0349f
C473 a_5960_42340# XA2.XA1.XA1.MN0.S 1.34e-19
C474 a_17408_41988# a_18560_41988# 0.00133f
C475 XA5.XA1.XA5.MN2.G EN 0.946f
C476 D<5> a_7328_44452# 1.48e-19
C477 XA8.XA7.MP0.G a_19928_44100# 2.31e-19
C478 XA2.XA1.XA5.MN2.G XA1.XA1.XA5.MP1.D 0.00329f
C479 XA0.XA7.MP0.G XA1.XA1.XA5.MN1.D 0.0102f
C480 XA3.XA4.MN0.G a_7328_47972# 0.155f
C481 D<1> a_18560_44804# 5.26e-19
C482 VREF a_9848_46564# 7.39e-19
C483 AVDD a_3440_40932# 0.00125f
C484 XA3.XA12.MP0.G a_8480_53252# 0.0661f
C485 XA4.XA11.MN1.G a_9848_53252# 0.0689f
C486 a_14888_53604# a_16040_53604# 0.00133f
C487 AVDD a_8480_52548# 0.00166f
C488 a_4808_40580# a_5960_40580# 0.00133f
C489 D<8> a_n232_45860# 0.162f
C490 XA5.XA1.XA5.MN2.G a_11000_41636# 0.0756f
C491 XA2.XA4.MN0.D XA2.XA1.XA5.MN0.D 9.9e-19
C492 CK_SAMPLE a_18560_50788# 0.157f
C493 XA4.XA10.MP0.G XA4.XA7.MP0.D 0.0601f
C494 XA20.XA4.MN0.D a_23600_52196# 0.056f
C495 XA4.XA9.MN1.G XA4.XA9.MN0.D 0.034f
C496 a_11000_52548# a_11000_52196# 0.0109f
C497 a_23600_52548# SARN 0.066f
C498 AVDD XA2.XA6.MN0.D 3.13e-19
C499 DONE a_21080_50436# 1.14e-19
C500 XB2.M1.G a_13808_1038# 0.00112f
C501 XB1.XA4.MP0.D a_8408_686# 0.0023f
C502 a_13808_1742# a_14960_1742# 0.00133f
C503 XB1.XA0.MP0.D a_9560_1390# 0.0719f
C504 XA20.XA3a.MN0.D a_22448_42692# 0.00125f
C505 a_13520_45508# EN 3.34e-19
C506 XA7.XA6.MP0.G a_14888_40580# 2.55e-19
C507 XA0.XA4.MN0.D XA0.XA1.XA1.MN0.D 0.00301f
C508 XA7.XA9.MN1.G XA7.XA6.MN0.D 0.0615f
C509 XA6.XA7.MP0.D a_14888_50436# 1.37e-19
C510 a_11000_51140# a_12368_51140# 8.89e-19
C511 XA3.XA1.XA5.MN2.G D<6> 0.624f
C512 AVDD a_9848_47268# 0.00125f
C513 XB1.XA4.MP0.D m3_7544_4532# 0.106f
C514 XB2.XA4.MP0.D XDAC2.XC1.XRES1A.B 0.377f
C515 EN XA3.XA1.XA4.MP1.D 0.0386f
C516 XA20.XA2a.MN0.D XA1.XA1.XA1.MN0.D 0.022f
C517 XA1.XA1.XA5.MN0.D a_2288_43396# 2.16e-19
C518 XA1.XA1.XA5.MP0.D a_3440_43396# 2.16e-19
C519 XA20.XA3.MN6.D XA20.XA3.MN1.D 0.159f
C520 AVDD a_23600_44100# 0.00154f
C521 a_5960_50436# VREF 0.0035f
C522 XA20.XA9.MP0.D a_23600_46212# 0.00334f
C523 XA1.XA6.MP0.D a_2288_49732# 0.00176f
C524 XA1.XA6.MP0.G a_3440_49732# 0.00239f
C525 D<8> li_14804_24912# 3.5e-20
C526 SARP a_9560_3150# 0.00116f
C527 XA4.XA1.XA4.MP0.D a_9848_42340# 2.16e-19
C528 XA4.XA1.XA4.MN0.D a_11000_42340# 2.16e-19
C529 EN a_5960_40228# 0.0674f
C530 D<1> a_17408_45860# 0.0774f
C531 XA5.XA1.XA5.MN2.G a_13520_45156# 1e-19
C532 XA6.XA1.XA5.MN2.G a_12368_45156# 0.00486f
C533 a_16040_48676# a_17408_48676# 8.89e-19
C534 XA6.XA6.MP0.G D<8> 0.0322f
C535 AVDD a_9848_41636# 0.00125f
C536 VREF a_7328_47620# 0.0671f
C537 XA2.XA4.MN0.D a_4808_47620# 0.0396f
C538 D<5> a_7328_45508# 0.00436f
C539 XA5.XA6.MP0.G XA3.XA3.MN0.G 0.0352f
C540 AVDD XA5.XA11.MP0.D 0.176f
C541 a_7328_53956# XA4.XA11.MN1.G 0.0295f
C542 XA8.XA1.XA1.MP2.D a_21080_40932# 0.00176f
C543 a_21080_41284# XA8.XA1.XA1.MP1.D 0.00176f
C544 a_9848_41284# a_9848_40932# 0.0109f
C545 D<2> a_14888_43044# 6.49e-19
C546 VREF a_21080_44452# 0.0179f
C547 XA20.XA3.MN0.D a_23600_44100# 0.0297f
C548 XA6.XA6.MP0.G a_14888_43748# 7.76e-20
C549 XA6.XA4.MN0.G a_16040_45860# 2.12e-19
C550 a_11000_46916# a_12368_46916# 8.89e-19
C551 D<6> XA2.XA1.XA4.MN1.D 0.00188f
C552 XA8.XA1.XA5.MN2.G a_17408_42692# 0.00442f
C553 XA7.XA1.XA5.MN2.G a_18560_42692# 0.0755f
C554 XA0.XA7.MP0.G XA0.XA1.XA4.MP0.D 0.00361f
C555 XA3.XA11.MN1.G XA3.XA8.MP0.D 6.42e-19
C556 XA2.XA10.MP0.D XA2.XA9.MN1.G 0.00406f
C557 XA7.XA11.MN1.G a_18560_51844# 3.12e-19
C558 a_9848_52900# a_9848_52548# 0.0109f
C559 AVDD D<7> 2.23f
C560 CK_SAMPLE XA0.XA7.MP0.G 0.0595f
C561 a_13808_3150# a_13808_2798# 0.0109f
C562 XA4.XA6.MP0.G a_9848_41284# 3.97e-20
C563 XA2.XA4.MN0.D a_4808_41988# 9.25e-20
C564 XA0.XA6.MP0.G XA0.XA1.XA1.MN0.D 0.00159f
C565 XA20.XA3a.MN0.D a_5960_43396# 0.00213f
C566 AVDD XDAC2.XC1.XRES1A.B 0.00509f
C567 XA5.XA1.XA5.MN2.D XA6.XA1.XA5.MN2.D 0.00869f
C568 a_13520_45508# a_13520_45156# 0.0109f
C569 CK_SAMPLE a_18560_49028# 7.31e-19
C570 AVDD a_8480_48324# 0.00131f
C571 a_21080_51844# a_21080_51492# 0.0109f
C572 SARN D<3> 0.027f
C573 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES16.B 0.0483f
C574 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES1A.B 0.00438f
C575 XDAC1.XC64b<1>.XRES8.B XDAC1.XC64b<1>.XRES2.B 0.44f
C576 XDAC2.XC64b<1>.XRES8.B li_14804_28392# 9.91e-20
C577 XA20.XA3a.MN0.D a_4808_40932# 0.0739f
C578 XA20.XA2a.MN0.D a_12368_41988# 0.00302f
C579 XA5.XA1.XA5.MN1.D a_12368_43748# 2.16e-19
C580 XA5.XA1.XA5.MP1.D a_13520_43748# 2.16e-19
C581 a_920_43748# a_2288_43748# 8.89e-19
C582 D<6> XDAC1.XC128b<2>.XRES16.B 3.2e-20
C583 XA0.XA6.MP2.G li_9184_19596# 3.5e-20
C584 EN XA0.XA1.XA5.MP0.D 0.0446f
C585 XA0.XA1.XA5.MP1.D XA0.XA1.XA2.MP0.D 6.52e-20
C586 XA0.XA1.XA5.MN1.D XA0.XA1.XA5.MN0.D 0.0488f
C587 a_13520_50788# XA5.XA6.MP0.G 1.75e-20
C588 AVDD a_12368_45156# 0.356f
C589 a_3440_50436# XA1.XA6.MP0.G 3.02e-20
C590 a_2288_50436# XA1.XA6.MP0.D 0.00176f
C591 a_920_51140# VREF 0.00383f
C592 XA6.XA1.XA5.MN2.G XA5.XA4.MN0.D 0.0939f
C593 SARN a_23600_48324# 0.0698f
C594 XA0.XA7.MP0.G a_920_49380# 0.00363f
C595 XDAC1.XC32a<0>.XRES8.B XDAC1.XC64a<0>.XRES8.B 6.7e-19
C596 XA1.XA4.MN0.D li_9184_9156# 0.00504f
C597 XA0.XA4.MN0.D XDAC1.XC1.XRES1B.B 0.00405f
C598 XA2.XA1.XA2.MP0.D a_5960_41636# 0.00224f
C599 XA6.XA1.XA2.MP0.D a_16040_41988# 0.0219f
C600 a_2288_42692# a_3440_42692# 0.00133f
C601 XA8.XA4.MN0.D a_21080_49028# 0.154f
C602 VREF a_5960_48676# 0.0191f
C603 a_9848_49380# a_9848_49028# 0.0109f
C604 D<7> a_2288_46564# 0.0695f
C605 XA5.XA1.XA5.MN2.G a_11000_46212# 0.00363f
C606 D<4> XA2.XA3.MN0.G 0.0259f
C607 AVDD a_19928_42692# 0.00159f
C608 AVDD a_18560_54308# 0.00166f
C609 a_920_54308# a_2288_54308# 8.89e-19
C610 SARP XDAC1.X16ab.XRES2.B 6.99f
C611 XA0.XA1.XA1.MN0.S a_920_41284# 0.0964f
C612 D<7> XA1.XA1.XA2.MP0.D 0.0132f
C613 a_4808_47620# a_4808_47268# 0.0109f
C614 XA6.XA4.MN0.G a_14888_46916# 0.0869f
C615 VREF a_21080_45508# 0.0556f
C616 AVDD a_16040_39876# 0.44f
C617 D<3> a_13520_43748# 6.49e-19
C618 a_21080_53252# a_22448_53252# 8.89e-19
C619 a_12368_53252# XA5.XA10.MP0.D 0.0677f
C620 AVDD a_11000_51844# 0.387f
C621 a_14888_53956# XA6.XA9.MN1.G 7.37e-20
C622 DONE XA8.XA7.MP0.D 0.217f
C623 XA2.XA11.MN1.G XA1.XA9.MN1.G 0.0169f
C624 D<5> a_8480_41284# 6.49e-19
C625 XA20.XA2a.MN0.D XA1.XA1.XA5.MN2.D 8.92e-20
C626 a_n232_45860# a_n232_45508# 0.0109f
C627 XA3.XA4.MN0.G a_8480_43748# 0.0157f
C628 XA20.XA3a.MN0.D EN 2.58f
C629 D<8> a_n232_44804# 0.043f
C630 XA7.XA3.MN0.G a_17408_45156# 0.0546f
C631 XA8.XA7.MP0.G XA8.XA1.XA1.MP1.D 0.144f
C632 XA3.XA1.XA5.MN2.G a_5960_40932# 0.0256f
C633 a_12368_52196# a_12368_51844# 0.0109f
C634 a_n232_52196# XA0.XA8.MP0.D 2.11e-19
C635 XA20.XA12.MP0.D VREF 0.00658f
C636 XA0.XA7.MP0.D a_n232_51844# 0.159f
C637 XA4.XA7.MP0.D XA5.XA7.MP0.D 0.00435f
C638 AVDD XA5.XA4.MN0.D 2.51f
C639 CK_SAMPLE a_18560_50084# 0.167f
C640 a_13808_n18# a_14960_n18# 0.00133f
C641 XA6.XA4.MN0.G XA6.XA1.XA1.MN0.S 5.22e-20
C642 a_12368_44452# EN 0.00173f
C643 a_18560_44452# a_18560_44100# 0.0109f
C644 XA20.XA2a.MN0.D XA8.XA1.XA4.MN1.D 0.00728f
C645 D<0> XA8.XA6.MN2.D 1.59e-19
C646 XA3.XA1.XA5.MN2.G XA3.XA6.MP0.G 0.0666f
C647 a_16040_51492# XA6.XA6.MP0.G 4.06e-20
C648 XA20.XA9.MP0.D a_21080_48324# 5.7e-20
C649 AVDD a_9848_46212# 0.00125f
C650 XA20.XA2a.MN0.D a_18560_40228# 2.1e-19
C651 a_18560_43396# a_18560_43044# 0.0109f
C652 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES1A.B 0.00405f
C653 XA20.XA9.MP0.D XA20.XA2.MN1.D 0.0349f
C654 XA1.XA6.MP0.G a_3440_48676# 0.0651f
C655 AVDD a_3440_43396# 0.00125f
C656 XA20.XA10.MN1.D a_23600_44100# 0.00405f
C657 XA5.XA6.MP0.G a_13520_49028# 0.0137f
C658 XA20.XA3.MN6.D a_22448_49380# 0.076f
C659 a_14888_49732# a_16040_49732# 0.00133f
C660 a_3440_49732# XA1.XA4.MN0.D 0.0659f
C661 SARP a_9560_334# 2.97e-20
C662 a_4808_41988# a_4808_41636# 0.0109f
C663 XA8.XA1.XA5.MN2.G a_19928_44100# 0.0709f
C664 XA4.XA1.XA5.MN2.G EN 0.897f
C665 XA8.XA4.MN0.D XA8.XA3.MN0.G 0.00642f
C666 XA0.XA7.MP0.G XA1.XA1.XA5.MP1.D 5.21e-20
C667 a_17408_48324# a_17408_47972# 0.0109f
C668 D<3> SARP 0.0407f
C669 D<1> a_17408_44804# 2.37e-19
C670 XA2.XA4.MN0.D a_5960_46564# 2.2e-19
C671 VREF a_8480_46564# 7.39e-19
C672 AVDD a_2288_40932# 0.358f
C673 a_2288_53604# XA1.XA11.MP0.D 0.00176f
C674 XA8.XA11.MN1.G XA8.XA11.MP0.D 0.0102f
C675 XA7.XA12.MP0.G XA7.XA11.MP0.D 0.0612f
C676 AVDD a_7328_52548# 0.405f
C677 XA3.XA12.MP0.G a_7328_53252# 0.00276f
C678 XA4.XA11.MN1.G a_8480_53252# 0.0238f
C679 a_17408_40932# a_17408_40580# 0.0109f
C680 XA6.XA3.MN0.G a_16040_46212# 0.155f
C681 XA6.XA4.MN0.G a_16040_44804# 5.54e-19
C682 XA5.XA1.XA5.MN2.G a_9848_41636# 0.128f
C683 XA2.XA4.MN0.D XA2.XA1.XA2.MP0.D 0.0111f
C684 VREF XA2.XA1.XA5.MP0.D 0.00202f
C685 XA0.XA11.MN1.G a_13808_2094# 0.00258f
C686 a_18560_46564# a_19928_46564# 8.89e-19
C687 a_5960_46564# a_5960_46212# 0.0109f
C688 CK_SAMPLE a_17408_50788# 0.00142f
C689 XA20.XA9.MP0.D a_23600_51844# 0.00348f
C690 XA20.XA4.MN0.D a_22448_52196# 2.16e-19
C691 AVDD XA2.XA6.MP0.G 5.93f
C692 DONE a_19928_50436# 6.41e-20
C693 XB2.M1.G a_12368_1038# 0.163f
C694 XB1.M1.G a_8408_686# 8.55e-20
C695 a_9560_1742# XB1.XA3.MN1.D 0.00176f
C696 XB1.XA0.MP0.D a_8408_1390# 0.0733f
C697 XB2.XA0.MP0.D XB2.XA3.MN1.D 0.193f
C698 XA20.XA3a.MN0.D a_21080_42692# 0.00156f
C699 XA20.XA2a.MN0.D XA4.XA1.XA2.MP0.D 0.223f
C700 a_12368_44804# a_13520_44804# 0.00133f
C701 a_n232_44804# a_n232_44452# 0.0109f
C702 XA2.XA4.MN0.G a_5960_42340# 1.28e-19
C703 XA3.XA1.XA5.MN2.D a_8480_44100# 0.0893f
C704 a_12368_45508# EN 1.42e-19
C705 XA7.XA6.MP0.G a_13520_40580# 1.4e-20
C706 SARN li_14804_24912# 0.00103f
C707 AVDD a_8480_47268# 0.00125f
C708 XA2.XA1.XA5.MN2.G D<6> 0.00595f
C709 XA7.XA9.MN1.G XA7.XA6.MP0.D 0.0618f
C710 a_17408_52900# VREF 0.00396f
C711 SARN XA6.XA6.MP0.G 0.0424f
C712 XB1.XA4.MP0.D m3_7472_4532# 0.0634f
C713 li_14804_23688# li_14804_23076# 0.00271f
C714 XDAC2.X16ab.XRES8.B XDAC2.XC128b<2>.XRES8.B 6.7e-19
C715 EN XA2.XA1.XA4.MP1.D 0.0386f
C716 XA20.XA2a.MN0.D XA1.XA1.XA1.MP1.D 0.00946f
C717 XA5.XA1.XA5.MP0.D XA5.XA1.XA5.MN0.D 0.00918f
C718 XA1.XA1.XA5.MP0.D a_2288_43396# 0.049f
C719 XA5.XA1.XA2.MP0.D XA6.XA1.XA2.MP0.D 0.00435f
C720 XA1.XA1.XA2.MP0.D a_3440_43396# 0.0961f
C721 a_16040_43748# a_16040_43396# 0.0109f
C722 SARN a_23600_47268# 0.0017f
C723 AVDD a_22448_44100# 0.37f
C724 XA5.XA6.MP0.G a_13520_50084# 6.4e-20
C725 XA5.XA6.MP0.D a_12368_50084# 0.049f
C726 XA1.XA6.MP0.G a_2288_49732# 0.099f
C727 XA20.XA3a.MN0.G XA20.XA3.MN1.D 0.0819f
C728 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES2.B 0.0136f
C729 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES8.B 0.471f
C730 XA3.XA3.MN0.G li_14804_25524# 0.00504f
C731 XA1.XA1.XA2.MP0.D a_2288_40932# 4.25e-20
C732 XA4.XA1.XA4.MN0.D a_9848_42340# 0.0474f
C733 a_22448_42692# a_22448_42340# 0.0109f
C734 XA6.XA1.XA5.MN2.G a_11000_45156# 7.1e-20
C735 XA5.XA1.XA5.MN2.G a_12368_45156# 7.1e-20
C736 a_3440_48676# a_3440_48324# 0.0109f
C737 AVDD a_8480_41636# 0.00125f
C738 VREF a_5960_47620# 0.0671f
C739 XA5.XA6.MP0.G XA2.XA3.MN0.G 0.0603f
C740 AVDD XA4.XA11.MP0.D 0.19f
C741 a_18560_53956# a_19928_53956# 8.89e-19
C742 a_8480_53956# XA3.XA11.MN1.G 0.00258f
C743 SARP li_9184_14472# 0.00103f
C744 XA3.XA1.XA1.MN0.S a_8480_40580# 0.00155f
C745 XA8.XA1.XA1.MN0.S a_21080_40932# 0.0271f
C746 VREF a_19928_44452# 7.12e-19
C747 SARN a_23600_41636# 5.16e-19
C748 XA6.XA4.MN0.G a_14888_45860# 0.0146f
C749 AVDD a_9560_1038# 0.00181f
C750 a_14888_47268# XA6.XA3.MN0.G 2.69e-19
C751 a_23600_47268# a_23600_46916# 0.0109f
C752 XA7.XA1.XA5.MN2.G a_17408_42692# 1.97e-19
C753 XA0.XA7.MP0.G XA0.XA1.XA4.MN0.D 7.2e-19
C754 XA7.XA11.MN1.G a_17408_51844# 4.48e-19
C755 a_21080_52900# XA8.XA10.MP0.G 0.0658f
C756 XA2.XA10.MP0.G XA3.XA10.MP0.G 0.00217f
C757 XA8.XA10.MP0.D a_21080_52548# 0.00224f
C758 AVDD XA0.XA6.MP2.D 0.172f
C759 CK_SAMPLE a_23600_51492# 7.93e-19
C760 a_8408_2798# a_9560_2798# 0.00133f
C761 XA4.XA4.MN0.G a_11000_43044# 0.0222f
C762 XA6.XA1.XA5.MN2.G a_14888_39876# 0.00169f
C763 XA20.XA3a.MN0.D a_4808_43396# 0.0736f
C764 AVDD XDAC1.XC1.XRES1A.B 0.00509f
C765 XA0.XA1.XA5.MN2.D a_920_45156# 0.155f
C766 XA4.XA7.MP0.D a_11000_51140# 0.00224f
C767 CK_SAMPLE a_17408_49028# 3.27e-19
C768 AVDD a_7328_48324# 0.359f
C769 XA4.XA8.MP0.D a_11000_51492# 0.00224f
C770 a_2288_51492# a_3440_51492# 0.00133f
C771 a_11000_51844# XA5.XA1.XA5.MN2.G 8.87e-19
C772 XA1.XA9.MN1.G a_3440_50788# 0.015f
C773 XA6.XA9.MN1.G XA6.XA6.MP2.D 0.0618f
C774 XA20.XA3a.MN0.D a_3440_40932# 0.0723f
C775 XA2.XA1.XA5.MN2.D a_5960_42692# 7.44e-20
C776 XA20.XA2a.MN0.D a_11000_41988# 0.00302f
C777 XA5.XA1.XA5.MP1.D a_12368_43748# 0.049f
C778 EN XA0.XA1.XA5.MN0.D 0.0063f
C779 XA0.XA1.XA5.MN1.D XA0.XA1.XA2.MP0.D 0.0102f
C780 a_12368_50788# XA5.XA6.MP0.G 1.34e-19
C781 a_14888_50436# a_16040_50436# 0.00133f
C782 AVDD a_11000_45156# 0.356f
C783 a_2288_50436# XA1.XA6.MP0.G 0.0678f
C784 XA0.XA6.MP2.G a_920_49732# 0.0109f
C785 XA5.XA1.XA5.MN2.G XA5.XA4.MN0.D 6.95e-19
C786 XA6.XA1.XA5.MN2.G XA4.XA4.MN0.D 6.95e-19
C787 XA0.XA1.XA4.MP1.D XA0.XA1.XA4.MP0.D 0.0488f
C788 XA2.XA1.XA2.MP0.D a_4808_41636# 0.00316f
C789 XA6.XA1.XA2.MP0.D a_14888_41988# 0.0568f
C790 XA5.XA1.XA4.MN1.D a_13520_42692# 0.0474f
C791 VREF a_4808_48676# 1.3e-19
C792 XA8.XA4.MN0.D a_19928_49028# 0.156f
C793 XA1.XA4.MN0.D a_3440_48676# 0.158f
C794 D<5> XA4.XA3.MN0.G 1.72e-19
C795 XA1.XA6.MP0.G a_3440_47620# 4.4e-19
C796 a_21080_49380# a_22448_49380# 8.89e-19
C797 D<4> XA1.XA3.MN0.G 0.0259f
C798 AVDD a_18560_42692# 0.00125f
C799 AVDD a_17408_54308# 0.448f
C800 XA4.XA1.XA1.MN0.S XA5.XA1.XA1.MN0.S 0.00217f
C801 XA0.XA1.XA1.MN0.S a_n232_41284# 0.0658f
C802 a_12368_41636# a_12368_41284# 0.0109f
C803 XA6.XA6.MP0.G SARP 0.0253f
C804 XA3.XA1.XA5.MN2.G a_5960_43396# 0.00442f
C805 a_16040_47620# a_17408_47620# 8.89e-19
C806 XA8.XA7.MP0.G XA8.XA1.XA5.MP0.D 0.00353f
C807 XA6.XA4.MN0.G a_13520_46916# 2.84e-19
C808 XA5.XA4.MN0.G a_14888_46916# 2.84e-19
C809 AVDD a_14888_39876# 0.00131f
C810 D<3> a_12368_43748# 7.77e-20
C811 XA4.XA11.MP0.D a_11000_52900# 0.00176f
C812 a_2288_53252# a_2288_52900# 0.0109f
C813 XA0.XA12.MP0.D XA1.XA9.MN0.D 1.35e-19
C814 AVDD a_9848_51844# 0.00166f
C815 a_11000_40228# a_11000_39876# 0.0109f
C816 D<5> a_7328_41284# 7.77e-20
C817 XA5.XA6.MP0.G a_13520_42340# 7.76e-20
C818 XA20.XA2a.MN0.D XA0.XA1.XA5.MN2.D 8.92e-20
C819 a_11000_45860# a_12368_45860# 8.89e-19
C820 XA1.XA6.MP0.G a_3440_41988# 7.76e-20
C821 XA3.XA4.MN0.G a_7328_43748# 6.3e-19
C822 XA8.XA7.MP0.G XA8.XA1.XA1.MN0.D 0.0378f
C823 XA3.XA1.XA5.MN2.G a_4808_40932# 6.44e-19
C824 XA8.XA1.XA5.MN2.G XA8.XA1.XA1.MP1.D 0.00107f
C825 XA2.XA1.XA5.MN2.G a_5960_40932# 1.69e-19
C826 XA6.XA9.MN1.G XA6.XA8.MP0.D 0.0132f
C827 AVDD XA4.XA4.MN0.D 2.51f
C828 CK_SAMPLE a_17408_50084# 0.00848f
C829 XA0.XA6.MP2.G li_9184_30036# 0.00508f
C830 D<6> XDAC1.XC0.XRES16.B 3.2e-20
C831 a_11000_44452# EN 0.00173f
C832 XA3.XA4.MN0.D a_8480_40228# 4.11e-20
C833 SARN XDAC2.XC32a<0>.XRES8.B 27.7f
C834 a_4808_44100# a_5960_44100# 0.00133f
C835 XA20.XA3a.MN0.D a_9848_41636# 0.00547f
C836 XA20.XA2a.MN0.D XA7.XA1.XA4.MN1.D 0.0128f
C837 XA4.XA6.MN2.D a_9848_50788# 0.0488f
C838 D<4> a_11000_50788# 0.161f
C839 XA0.XA6.MN2.D a_n232_50436# 0.00176f
C840 a_920_51140# XA0.XA6.MP0.G 6.76e-20
C841 XA0.XA6.MP2.G a_920_50436# 0.0879f
C842 AVDD a_8480_46212# 0.00125f
C843 XA6.XA9.MN1.G a_16040_49380# 2.54e-19
C844 li_9184_18564# li_9184_17952# 0.00271f
C845 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES2.B 0.0307f
C846 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES16.B 0.0381f
C847 XDAC1.XC128b<2>.XRES1A.B XDAC1.XC128a<1>.XRES1A.B 0.00444f
C848 SARP a_23600_41636# 0.161f
C849 XA7.XA1.XA2.MP0.D XA7.XA1.XA4.MN1.D 0.056f
C850 a_4808_43044# a_5960_43044# 0.00133f
C851 XA0.XA6.MP0.G li_14804_9156# 1.85e-20
C852 EN a_22448_42340# 5.7e-20
C853 XA1.XA6.MP0.G a_2288_48676# 0.0881f
C854 D<0> XA8.XA4.MN0.G 0.239f
C855 D<7> XA20.XA3a.MN0.D 0.0703f
C856 XA20.XA9.MP0.D a_23600_45156# 0.00558f
C857 AVDD a_2288_43396# 0.361f
C858 XA20.XA10.MN1.D a_22448_44100# 1.87e-19
C859 SARN a_23600_46212# 0.0017f
C860 XA5.XA6.MP0.G a_12368_49028# 0.0307f
C861 a_19928_50084# XA8.XA4.MN0.D 3.12e-20
C862 XA20.XA3a.MN0.G a_22448_49380# 0.0948f
C863 a_2288_49732# XA1.XA4.MN0.D 0.0674f
C864 a_16040_41988# a_17408_41988# 8.89e-19
C865 XA8.XA1.XA5.MN2.G a_18560_44100# 2.31e-19
C866 XA3.XA1.XA5.MN2.G EN 0.946f
C867 XA0.XA7.MP0.G XA0.XA1.XA5.MP1.D 0.00329f
C868 XA2.XA4.MN0.G a_5960_47972# 0.155f
C869 VREF a_7328_46564# 0.0175f
C870 XA2.XA4.MN0.D a_4808_46564# 0.001f
C871 AVDD a_920_40932# 0.358f
C872 a_13520_53604# a_14888_53604# 8.89e-19
C873 XA8.XA11.MN1.G XA7.XA11.MP0.D 0.0114f
C874 AVDD a_5960_52548# 0.405f
C875 XA4.XA11.MN1.G a_7328_53252# 3.16e-19
C876 XA3.XA11.MN1.G a_9848_53252# 2.81e-19
C877 a_3440_40580# a_4808_40580# 8.89e-19
C878 XA6.XA3.MN0.G a_14888_46212# 0.157f
C879 XA6.XA4.MN0.G a_14888_44804# 0.00858f
C880 XA4.XA1.XA5.MN2.G a_9848_41636# 0.00417f
C881 XA0.XA11.MN1.G a_12368_2094# 0.156f
C882 AVDD XA1.XA6.MN0.D 3.13e-19
C883 CK_SAMPLE a_16040_50788# 0.00142f
C884 XA3.XA10.MP0.G XA3.XA7.MP0.D 0.0601f
C885 a_9848_52548# a_9848_52196# 0.0109f
C886 a_9560_1742# XB1.XA3.MN0.S 0.0687f
C887 a_12368_1742# a_13808_1742# 8e-19
C888 XB2.XA0.MP0.D XB2.XA3.MN0.S 0.572f
C889 a_8408_1742# XB1.XA3.MN1.D 0.00685f
C890 SAR_IP a_11000_334# 0.0566f
C891 XA20.XA3a.MN0.D a_19928_42692# 0.00778f
C892 XA2.XA6.MP0.G a_5960_40228# 5.5e-19
C893 XA6.XA6.MP0.G a_16040_40580# 5.5e-19
C894 XA2.XA4.MN0.G a_4808_42340# 7.97e-19
C895 XA3.XA1.XA5.MN2.D a_7328_44100# 0.124f
C896 a_11000_45508# EN 1.42e-19
C897 XA7.XA6.MP0.G a_12368_40580# 1.86e-20
C898 XA8.XA7.MP0.G a_22448_51140# 0.00105f
C899 a_9848_51140# a_11000_51140# 0.00133f
C900 AVDD a_7328_47268# 0.356f
C901 XA2.XA1.XA5.MN2.G XA1.XA6.MN2.D 6.33e-19
C902 XA0.XA7.MP0.G D<6> 4.48e-21
C903 a_16040_52900# VREF 0.00396f
C904 XA7.XA9.MN1.G XA7.XA6.MP0.G 0.0725f
C905 XA1.XA9.MN1.G a_3440_50084# 0.00969f
C906 XA5.XA7.MP0.D a_13520_50436# 1.37e-19
C907 EN XA2.XA1.XA4.MN1.D 3.17e-19
C908 XA20.XA2a.MN0.D XA0.XA1.XA1.MP1.D 0.00946f
C909 XA5.XA1.XA2.MP0.D XA5.XA1.XA5.MN0.D 0.056f
C910 AVDD a_21080_44100# 0.359f
C911 D<0> a_21080_49380# 0.00891f
C912 XA5.XA6.MP0.G a_12368_50084# 0.159f
C913 XA0.XA6.MP2.G a_920_48676# 0.00918f
C914 D<4> a_11000_49028# 0.00884f
C915 XA20.XA3a.MN0.G XA20.XA3.MN6.D 1.76f
C916 D<8> XDAC2.X16ab.XRES8.B 4.06e-21
C917 SARP XB1.XA2.MN0.G 0.00236f
C918 XA5.XA1.XA5.MN2.G a_11000_45156# 0.00486f
C919 XA8.XA4.MN0.D a_21080_47972# 0.0546f
C920 a_14888_48676# a_16040_48676# 0.00133f
C921 AVDD a_7328_41636# 0.404f
C922 XA4.XA6.MP0.G XA4.XA3.MN0.G 0.0501f
C923 XA7.XA6.MP0.G a_18560_46916# 5e-19
C924 XA1.XA4.MN0.D a_3440_47620# 0.0396f
C925 VREF a_4808_47620# 7.12e-19
C926 XA5.XA6.MP0.G XA1.XA3.MN0.G 0.0267f
C927 AVDD XA3.XA11.MP0.D 0.176f
C928 a_5960_53956# XA2.XA12.MP0.G 0.0658f
C929 a_7328_53956# XA3.XA11.MN1.G 0.00198f
C930 XA20.XA12.MP0.D a_23600_53604# 0.0674f
C931 XA3.XA1.XA1.MN0.S a_7328_40580# 0.0318f
C932 a_19928_41284# XA8.XA1.XA1.MN0.D 0.00224f
C933 a_8480_41284# a_8480_40932# 0.0109f
C934 VREF a_18560_44452# 7.12e-19
C935 XA1.XA6.MP0.G XA1.XA1.XA5.MN0.D 7.41e-19
C936 XA5.XA4.MN0.G a_14888_45860# 2.2e-19
C937 XA6.XA4.MN0.G a_13520_45860# 2.2e-19
C938 AVDD a_8408_1038# 0.488f
C939 a_9848_46916# a_11000_46916# 0.00133f
C940 XA7.XA1.XA5.MN2.G a_16040_42692# 0.00442f
C941 XA7.XA11.MN1.G a_16040_51844# 2.62e-19
C942 a_8480_52900# a_8480_52548# 0.0109f
C943 a_19928_52900# XA8.XA10.MP0.G 0.0681f
C944 XA8.XA10.MP0.D a_19928_52548# 0.00316f
C945 a_14888_53252# XA6.XA9.MN1.G 5.25e-19
C946 AVDD XA0.XA6.MN2.D 3.77e-19
C947 CK_SAMPLE a_22448_51492# 0.00729f
C948 XA4.XA4.MN0.G a_9848_43044# 0.0409f
C949 XA20.XA2a.MN0.D a_23600_44452# 0.0026f
C950 XA6.XA1.XA5.MN2.G a_13520_39876# 2.97e-20
C951 SARN CK_SAMPLE_BSSW 0.00161f
C952 XA1.XA4.MN0.D a_3440_41988# 9.24e-20
C953 XA8.XA3.MN0.G EN 0.00979f
C954 XA20.XA3a.MN0.D a_3440_43396# 0.0723f
C955 XA4.XA1.XA5.MN2.D XA5.XA1.XA5.MN2.D 0.00869f
C956 XA0.XA1.XA5.MN2.D a_n232_45156# 0.153f
C957 a_12368_45508# a_12368_45156# 0.0109f
C958 XA1.XA9.MN1.G a_2288_50788# 0.00281f
C959 XA4.XA7.MP0.D a_9848_51140# 0.00388f
C960 CK_SAMPLE a_16040_49028# 3.27e-19
C961 AVDD a_5960_48324# 0.359f
C962 XA4.XA8.MP0.D a_9848_51492# 0.00224f
C963 a_19928_51844# a_19928_51492# 0.0109f
C964 XA6.XA9.MN1.G XA6.XA6.MN2.D 0.126f
C965 a_2288_53604# VREF 0.00396f
C966 li_14804_29004# li_14804_28392# 0.00271f
C967 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES2.B 0.0307f
C968 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES16.B 0.0381f
C969 XDAC2.XC0.XRES1A.B XDAC2.XC64b<1>.XRES1A.B 0.00444f
C970 XDAC1.XC64b<1>.XRES8.B li_9184_28392# 9.91e-20
C971 XA20.XA3a.MN0.D a_2288_40932# 0.0674f
C972 XA20.XA2a.MN0.D a_9848_41988# 0.0844f
C973 a_n232_43748# a_920_43748# 0.00133f
C974 XA0.XA6.MP2.G XDAC1.XC128b<2>.XRES1A.B 4.06e-21
C975 a_19928_44452# XA8.XA1.XA2.MP0.D 5.16e-20
C976 a_9848_44100# XA4.XA1.XA2.MP0.D 2.92e-19
C977 EN XA0.XA1.XA2.MP0.D 0.156f
C978 AVDD a_9848_45156# 0.00125f
C979 XA8.XA7.MP0.G VREF 0.687f
C980 XA0.XA6.MP2.G a_n232_49732# 7.01e-19
C981 XA5.XA1.XA5.MN2.G XA4.XA4.MN0.D 0.0939f
C982 D<4> a_11000_50084# 0.0155f
C983 li_9184_13248# li_9184_12636# 0.00271f
C984 EN a_12368_41284# 0.00564f
C985 XA1.XA4.MN0.D XDAC1.XC64a<0>.XRES1A.B 0.00405f
C986 XA0.XA4.MN0.D li_9184_9156# 1.85e-20
C987 XA5.XA1.XA4.MN1.D a_12368_42692# 2.16e-19
C988 XA5.XA1.XA4.MP1.D a_13520_42692# 2.16e-19
C989 a_920_42692# a_2288_42692# 8.89e-19
C990 XA20.XA3a.MN0.G XA8.XA4.MN0.G 0.00652f
C991 D<5> XA3.XA3.MN0.G 1.2f
C992 XA1.XA6.MP0.G a_2288_47620# 6.35e-19
C993 a_8480_49380# a_8480_49028# 0.0109f
C994 D<4> D<8> 0.0323f
C995 AVDD a_17408_42692# 0.358f
C996 XA2.XA6.MP0.G XA20.XA3a.MN0.D 0.0687f
C997 XA5.XA6.MP0.G a_13520_47972# 6.28e-19
C998 XA1.XA4.MN0.D a_2288_48676# 0.154f
C999 VREF a_3440_48676# 1.3e-19
C1000 a_n232_54308# a_920_54308# 0.00133f
C1001 AVDD a_16040_54308# 0.447f
C1002 SARP li_9184_24912# 0.00103f
C1003 XA4.XA1.XA1.MN0.S XA4.XA1.XA1.MP2.D 0.0708f
C1004 XA3.XA1.XA5.MN2.G a_4808_43396# 1.95e-19
C1005 a_3440_47620# a_3440_47268# 0.0109f
C1006 XA8.XA7.MP0.G XA8.XA1.XA5.MN0.D 7.2e-19
C1007 XA5.XA4.MN0.G a_13520_46916# 0.0885f
C1008 AVDD a_13520_39876# 0.00131f
C1009 XA3.XA6.MP0.G a_8480_44452# 7.76e-20
C1010 AVDD a_8480_51844# 0.00166f
C1011 XA0.XA12.MP0.D XA1.XA9.MN1.G 0.00349f
C1012 a_19928_53252# a_21080_53252# 0.00133f
C1013 a_11000_53252# XA4.XA10.MP0.D 0.0661f
C1014 XA6.XA11.MN1.G a_14888_52548# 2.85e-19
C1015 a_22448_40228# a_23600_40228# 0.00133f
C1016 XA5.XA6.MP0.G a_12368_42340# 5.5e-19
C1017 XA20.XA2a.MN0.D a_23600_45508# 0.0688f
C1018 a_23600_46212# a_23600_45860# 0.0109f
C1019 XA1.XA6.MP0.G a_2288_41988# 5.5e-19
C1020 XA20.XA3a.MN0.D a_22448_44100# 0.00697f
C1021 XA6.XA3.MN0.G a_16040_45156# 0.0546f
C1022 XA8.XA1.XA5.MN2.G XA8.XA1.XA1.MN0.D 0.0288f
C1023 XA2.XA1.XA5.MN2.G a_4808_40932# 0.00729f
C1024 XA3.XA4.MN0.D XA3.XA1.XA4.MN1.D 9.89e-19
C1025 SARN a_23600_51844# 0.156f
C1026 a_11000_52196# a_11000_51844# 0.0109f
C1027 XA2.XA9.MN1.G a_5960_51492# 6.57e-19
C1028 a_22448_55012# VREF 0.0015f
C1029 a_7328_52548# XA4.XA1.XA5.MN2.G 1.75e-19
C1030 XA3.XA7.MP0.D XA4.XA7.MP0.D 0.00435f
C1031 AVDD XA3.XA4.MN0.D 2.65f
C1032 CK_SAMPLE a_16040_50084# 0.00848f
C1033 a_12368_n18# a_13808_n18# 8e-19
C1034 a_9848_44452# EN 0.00154f
C1035 XA3.XA4.MN0.D a_7328_40228# 4.07e-20
C1036 a_17408_44452# a_17408_44100# 0.0109f
C1037 XA20.XA3a.MN0.D a_8480_41636# 0.00547f
C1038 XA20.XA2a.MN0.D XA7.XA1.XA4.MP1.D 0.0128f
C1039 XA5.XA1.XA5.MN2.D XA5.XA1.XA2.MP0.D 4.72e-19
C1040 XA0.XA6.MP2.G a_n232_50436# 5.7e-19
C1041 a_17408_52196# VREF 0.00396f
C1042 XA4.XA1.XA5.MN2.G XA2.XA6.MP0.G 3.47e-19
C1043 AVDD a_7328_46212# 0.356f
C1044 XA6.XA9.MN1.G a_14888_49380# 4.23e-20
C1045 XA7.XA1.XA2.MP0.D XA7.XA1.XA4.MP1.D 4.34e-19
C1046 a_17408_43396# a_17408_43044# 0.0109f
C1047 EN a_21080_42340# 0.159f
C1048 XA1.XA6.MP0.G li_14804_9768# 0.00504f
C1049 XA0.XA6.MP2.G a_920_47620# 0.0147f
C1050 AVDD a_920_43396# 0.361f
C1051 a_13520_49732# a_14888_49732# 8.89e-19
C1052 a_2288_49732# VREF 0.029f
C1053 SARP CK_SAMPLE_BSSW 0.00161f
C1054 a_3440_41988# a_3440_41636# 0.0109f
C1055 XA8.XA1.XA5.MN2.G a_17408_44100# 0.00556f
C1056 XA7.XA1.XA5.MN2.G a_18560_44100# 0.0693f
C1057 a_16040_48324# a_16040_47972# 0.0109f
C1058 XA2.XA4.MN0.G a_4808_47972# 0.153f
C1059 XA0.XA7.MP0.G XA0.XA1.XA5.MN1.D 6.68e-19
C1060 XA2.XA1.XA5.MN2.G EN 0.897f
C1061 XA3.XA6.MP0.G a_8480_45508# 7.76e-20
C1062 XA7.XA4.MN0.G XA8.XA4.MN0.G 0.12f
C1063 XA7.XA6.MP0.G a_18560_45860# 1.38e-19
C1064 VREF a_5960_46564# 0.0175f
C1065 AVDD a_n232_40932# 0.00125f
C1066 XA7.XA4.MN0.D XA7.XA3.MN0.G 0.00642f
C1067 XA20.XA12.MP0.G XA8.XA10.MP0.G 9.09e-19
C1068 a_920_53604# XA0.XA11.MP0.D 0.00176f
C1069 AVDD a_4808_52548# 0.00166f
C1070 XA3.XA11.MN1.G a_8480_53252# 0.0758f
C1071 XA6.XA1.XA1.MN0.D a_14888_40228# 0.00155f
C1072 a_16040_40932# a_16040_40580# 0.0109f
C1073 XA6.XA4.MN0.G a_13520_44804# 2.2e-19
C1074 XA5.XA4.MN0.G a_14888_44804# 2.2e-19
C1075 D<4> a_11000_42340# 7.76e-20
C1076 XA4.XA1.XA5.MN2.G a_8480_41636# 0.131f
C1077 XA0.XA6.MP2.G a_920_41988# 7.76e-20
C1078 XA1.XA4.MN0.D XA1.XA1.XA5.MN0.D 9.89e-19
C1079 XA0.XA11.MN1.G a_11000_2094# 0.156f
C1080 XA2.XA6.MP0.G XA2.XA1.XA4.MP1.D 0.00121f
C1081 a_17408_46564# a_18560_46564# 0.00133f
C1082 a_4808_46564# a_4808_46212# 0.0109f
C1083 XA6.XA6.MP0.G a_16040_43044# 5.5e-19
C1084 CK_SAMPLE a_14888_50788# 0.157f
C1085 XA8.XA10.MP0.G a_21080_52196# 0.0441f
C1086 XA3.XA9.MN1.G XA4.XA9.MN1.G 0.0531f
C1087 AVDD XA1.XA6.MP0.D 0.144f
C1088 XB2.XA4.MP0.D a_14960_1390# 0.00559f
C1089 a_14960_2094# XB2.XA3.MN1.D 0.00291f
C1090 SAR_IN CK_SAMPLE_BSSW 0.0123f
C1091 SAR_IP a_9560_334# 1.73e-19
C1092 XA20.XA3a.MN0.D a_18560_42692# 0.01f
C1093 XA2.XA6.MP0.G a_4808_40228# 7.76e-20
C1094 XA20.XA2.MN1.D SARP 0.11f
C1095 a_11000_44804# a_12368_44804# 8.89e-19
C1096 XA6.XA6.MP0.G a_14888_40580# 7.76e-20
C1097 XA8.XA4.MN0.G XA8.XA1.XA4.MN0.D 0.00331f
C1098 XA4.XA3.MN0.G a_9848_43396# 6.8e-20
C1099 a_9848_45508# EN 3.34e-19
C1100 SARN XDAC2.X16ab.XRES8.B 27.7f
C1101 a_12368_51492# D<3> 2.41e-19
C1102 XA8.XA7.MP0.G a_21080_51140# 0.077f
C1103 AVDD a_5960_47268# 0.356f
C1104 XA2.XA1.XA5.MN2.G XA1.XA6.MP2.D 0.00313f
C1105 XA1.XA9.MN1.G a_2288_50084# 0.00281f
C1106 li_9184_23688# li_9184_23076# 0.00271f
C1107 XDAC1.X16ab.XRES8.B XDAC1.XC128b<2>.XRES8.B 6.7e-19
C1108 XA3.XA3.MN0.G a_9848_40932# 9.08e-19
C1109 XA0.XA6.MP0.G li_14804_19596# 0.00504f
C1110 EN XA1.XA1.XA4.MN1.D 3.17e-19
C1111 XA20.XA2a.MN0.D XA0.XA1.XA1.MN0.D 0.0221f
C1112 XA5.XA1.XA2.MP0.D XA5.XA1.XA5.MP0.D 4.34e-19
C1113 a_14888_43748# a_14888_43396# 0.0109f
C1114 AVDD a_19928_44100# 0.00159f
C1115 a_2288_50436# VREF 0.0035f
C1116 D<0> a_19928_49380# 5.91e-19
C1117 XA0.XA6.MP2.G a_n232_48676# 3.48e-19
C1118 XA4.XA1.XA5.MN2.G a_7328_48324# 0.00455f
C1119 D<4> a_9848_49028# 5.7e-19
C1120 XA0.XA6.MP0.D a_920_49732# 0.00176f
C1121 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES2.B 0.0136f
C1122 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES8.B 0.471f
C1123 XA3.XA3.MN0.G XDAC2.X16ab.XRES4.B 0.00405f
C1124 SARP a_9560_3502# 0.00116f
C1125 XA8.XA1.XA2.MP0.D a_21080_41284# 1.07e-19
C1126 XA8.XA1.XA4.MN0.D XA8.XA1.XA4.MP0.D 0.00918f
C1127 a_7328_43044# XA3.XA1.XA1.MN0.S 4.06e-20
C1128 XA3.XA1.XA4.MN0.D a_8480_42340# 0.0474f
C1129 a_21080_42692# a_21080_42340# 0.0109f
C1130 EN a_2288_40228# 0.0658f
C1131 XA5.XA1.XA5.MN2.G a_9848_45156# 1.95e-19
C1132 XA8.XA4.MN0.D a_19928_47972# 0.0788f
C1133 a_2288_48676# a_2288_48324# 0.0109f
C1134 AVDD a_5960_41636# 0.404f
C1135 XA4.XA6.MP0.G XA3.XA3.MN0.G 0.271f
C1136 XA7.XA6.MP0.G a_17408_46916# 5.5e-19
C1137 XA1.XA4.MN0.D a_2288_47620# 0.00498f
C1138 VREF a_3440_47620# 7.12e-19
C1139 XA5.XA6.MP0.G D<8> 0.033f
C1140 XA1.XA6.MP0.G a_3440_46564# 7.76e-20
C1141 a_19928_54308# XA8.XA11.MN1.G 2.9e-19
C1142 AVDD XA2.XA11.MP0.D 0.19f
C1143 a_17408_53956# a_18560_53956# 0.00133f
C1144 a_4808_53956# XA2.XA12.MP0.G 0.0704f
C1145 a_5960_53956# XA3.XA11.MN1.G 0.0442f
C1146 XA20.XA12.MP0.D a_22448_53604# 0.0694f
C1147 XA20.XA12.MP0.G a_21080_53604# 0.00586f
C1148 SARP XDAC1.XC32a<0>.XRES8.B 27.7f
C1149 VREF a_17408_44452# 0.0182f
C1150 XA1.XA6.MP0.G XA1.XA1.XA5.MP0.D 0.00121f
C1151 XA5.XA4.MN0.G a_13520_45860# 0.0146f
C1152 AVDD a_14960_1390# 0.434f
C1153 a_13520_47268# XA5.XA3.MN0.G 2.69e-19
C1154 a_22448_47268# a_22448_46916# 0.0109f
C1155 XA6.XA1.XA5.MN2.G a_16040_42692# 1.97e-19
C1156 XA7.XA1.XA5.MN2.G a_14888_42692# 1.95e-19
C1157 XA1.XA10.MP0.D XA1.XA9.MN1.G 0.00406f
C1158 XA1.XA10.MP0.G XA2.XA10.MP0.G 0.00217f
C1159 AVDD XA0.XA6.MP2.G 2.23f
C1160 CK_SAMPLE a_21080_51492# 0.00287f
C1161 XA7.XA6.MP0.G XA7.XA1.XA1.MN0.S 0.0145f
C1162 XA20.XA2a.MN0.D a_22448_44452# 0.00148f
C1163 XA5.XA1.XA5.MN2.G a_13520_39876# 0.00325f
C1164 XA6.XA1.XA5.MN2.G a_12368_39876# 8.8e-19
C1165 D<7> a_3440_40228# 2.88e-19
C1166 XA1.XA4.MN0.D a_2288_41988# 9.15e-20
C1167 XA7.XA3.MN0.G EN 0.00979f
C1168 XA2.XA3.MN0.G XA2.XA1.XA5.MN1.D 8.47e-19
C1169 XA20.XA3a.MN0.D a_2288_43396# 0.00213f
C1170 D<3> a_13520_40580# 5.26e-19
C1171 CK_SAMPLE a_14888_49028# 7.31e-19
C1172 AVDD a_4808_48324# 0.00131f
C1173 a_920_51492# a_2288_51492# 8.89e-19
C1174 a_5960_52196# D<6> 7.56e-20
C1175 SARN D<4> 0.027f
C1176 XA6.XA9.MN1.G D<2> 0.0378f
C1177 a_920_53604# VREF 0.00351f
C1178 XA20.XA3a.MN0.D a_920_40932# 0.0658f
C1179 XA20.XA2a.MN0.D a_8480_41988# 0.0861f
C1180 XA4.XA1.XA5.MP1.D a_11000_43748# 0.049f
C1181 a_13520_50436# a_14888_50436# 8.89e-19
C1182 AVDD a_8480_45156# 0.00125f
C1183 a_920_50436# XA0.XA6.MP0.D 0.00176f
C1184 XA8.XA1.XA5.MN2.G VREF 0.704f
C1185 D<4> a_9848_50084# 5.7e-19
C1186 D<0> XA8.XA6.MP0.D 0.0323f
C1187 EN a_11000_41284# 0.00564f
C1188 XA0.XA1.XA4.MN1.D XA0.XA1.XA4.MN0.D 0.0488f
C1189 XA5.XA1.XA4.MP1.D a_12368_42692# 0.049f
C1190 SARN a_23600_45156# 0.00206f
C1191 D<2> a_16040_46916# 0.0185f
C1192 D<5> XA2.XA3.MN0.G 0.026f
C1193 a_19928_49380# a_21080_49380# 0.00133f
C1194 AVDD a_16040_42692# 0.358f
C1195 XA5.XA6.MP0.G a_12368_47972# 8.92e-19
C1196 VREF a_2288_48676# 0.0191f
C1197 XA7.XA4.MN0.D a_18560_49028# 0.156f
C1198 AVDD a_14888_54308# 0.00166f
C1199 a_11000_41636# a_11000_41284# 0.0109f
C1200 VREF a_17408_45508# 0.0556f
C1201 XA7.XA6.MP0.G a_18560_44804# 7.76e-20
C1202 XA2.XA1.XA5.MN2.G a_4808_43396# 0.00504f
C1203 a_14888_47620# a_16040_47620# 0.00133f
C1204 XA8.XA7.MP0.G XA8.XA1.XA2.MP0.D 0.144f
C1205 XA5.XA4.MN0.G a_12368_46916# 0.0662f
C1206 AVDD a_12368_39876# 0.438f
C1207 XA3.XA6.MP0.G a_7328_44452# 5.5e-19
C1208 AVDD a_7328_51844# 0.387f
C1209 XA0.XA12.MP0.G XA0.XA9.MN1.G 4.5e-19
C1210 a_9848_53252# XA4.XA10.MP0.D 0.0692f
C1211 a_920_53252# a_920_52900# 0.0109f
C1212 XA6.XA11.MN1.G a_13520_52548# 9.76e-19
C1213 a_9848_40228# a_9848_39876# 0.0109f
C1214 XA20.XA2a.MN0.D a_22448_45508# 0.0445f
C1215 a_9848_45860# a_11000_45860# 0.00133f
C1216 XA2.XA4.MN0.G a_5960_43748# 6.3e-19
C1217 XA8.XA4.MN0.G XA8.XA1.XA5.MP1.D 0.00138f
C1218 XA6.XA3.MN0.G a_14888_45156# 0.0805f
C1219 XA20.XA3a.MN0.D a_21080_44100# 6.57e-19
C1220 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.D 0.0825f
C1221 XA2.XA1.XA5.MN2.G a_3440_40932# 0.00838f
C1222 XA3.XA4.MN0.D XA3.XA1.XA4.MP1.D 9.71e-19
C1223 AVDD XA2.XA4.MN0.D 2.65f
C1224 CK_SAMPLE a_14888_50084# 0.167f
C1225 XA2.XA9.MN1.G a_4808_51492# 0.0118f
C1226 XA5.XA4.MN0.G XA5.XA1.XA1.MN0.S 5.22e-20
C1227 XA0.XA6.MP2.G XDAC1.XC0.XRES1A.B 0.00406f
C1228 a_8480_44452# EN 0.00154f
C1229 a_3440_44100# a_4808_44100# 8.89e-19
C1230 SARN li_14804_15084# 0.00103f
C1231 XA20.XA2a.MN0.D XA6.XA1.XA4.MP1.D 0.0128f
C1232 a_4808_45156# XA2.XA1.XA2.MP0.D 1.56e-20
C1233 a_16040_52196# VREF 0.00396f
C1234 XA3.XA1.XA5.MN2.G XA2.XA6.MP0.G 0.093f
C1235 AVDD a_5960_46212# 0.356f
C1236 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES8.B 0.471f
C1237 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES2.B 0.0136f
C1238 XA20.XA2a.MN0.D a_14888_40228# 2.1e-19
C1239 XA3.XA1.XA2.MP0.D a_8480_42692# 0.0946f
C1240 a_3440_43044# a_4808_43044# 8.89e-19
C1241 XA0.XA6.MP0.G XDAC2.XC64a<0>.XRES1A.B 2.23e-21
C1242 XA0.XA4.MN0.D li_9184_19596# 0.00504f
C1243 XA4.XA1.XA5.MN2.G a_7328_47268# 0.00363f
C1244 AVDD a_n232_43396# 0.00125f
C1245 a_18560_50084# XA7.XA4.MN0.D 3.12e-20
C1246 a_920_49732# VREF 0.029f
C1247 XA0.XA6.MP2.G a_n232_47620# 5.21e-19
C1248 D<4> a_11000_47972# 0.0147f
C1249 a_14888_41988# a_16040_41988# 0.00133f
C1250 XA0.XA7.MP0.G EN 0.963f
C1251 XA8.XA1.XA5.MN2.G a_16040_44100# 7.1e-20
C1252 XA7.XA1.XA5.MN2.G a_17408_44100# 7.1e-20
C1253 XA3.XA6.MP0.G a_7328_45508# 5.5e-19
C1254 D<6> a_5960_44452# 1.47e-19
C1255 D<4> SARP 0.0406f
C1256 XA7.XA6.MP0.G a_17408_45860# 5.5e-19
C1257 XA1.XA4.MN0.D a_3440_46564# 0.001f
C1258 VREF a_4808_46564# 7.39e-19
C1259 AVDD XA8.XA1.XA1.MP1.D 0.0604f
C1260 a_12368_53604# a_13520_53604# 0.00133f
C1261 a_920_53604# XA0.XA11.MN1.G 0.0658f
C1262 XA6.XA12.MP0.G XA6.XA11.MP0.D 0.0612f
C1263 XA7.XA11.MN1.G XA7.XA11.MP0.D 0.0383f
C1264 AVDD a_3440_52548# 0.00166f
C1265 XA3.XA11.MN1.G a_7328_53252# 0.0762f
C1266 XA2.XA12.MP0.G a_5960_53252# 0.00276f
C1267 a_2288_40580# a_3440_40580# 0.00133f
C1268 XA5.XA3.MN0.G a_13520_46212# 0.157f
C1269 XA1.XA4.MN0.D XA1.XA1.XA5.MP0.D 9.71e-19
C1270 D<4> a_9848_42340# 6.49e-19
C1271 XA4.XA1.XA5.MN2.G a_7328_41636# 0.0736f
C1272 XA3.XA1.XA5.MN2.G a_8480_41636# 0.0039f
C1273 XA0.XA6.MP2.G a_n232_41988# 6.49e-19
C1274 XA0.XA11.MN1.G a_9560_2094# 0.00258f
C1275 XA2.XA6.MP0.G XA2.XA1.XA4.MN1.D 7.41e-19
C1276 XA6.XA6.MP0.G a_14888_43044# 7.76e-20
C1277 XA5.XA4.MN0.G a_13520_44804# 0.00858f
C1278 CK_SAMPLE a_13520_50788# 0.157f
C1279 XA2.XA10.MP0.G XA2.XA7.MP0.D 0.0601f
C1280 XA8.XA10.MP0.G a_19928_52196# 0.0131f
C1281 a_8480_52548# a_8480_52196# 0.0109f
C1282 a_19928_52548# XA8.XA9.MN0.D 0.00176f
C1283 a_21080_52548# XA8.XA9.MN1.G 0.0658f
C1284 XA3.XA9.MN1.G XA3.XA9.MN0.D 0.034f
C1285 AVDD XA1.XA6.MP0.G 5.92f
C1286 a_11000_1742# a_12368_1742# 8.89e-19
C1287 XB1.XA0.MP0.D XB1.XA3.MN1.D 0.193f
C1288 XA20.XA3a.MN0.D a_17408_42692# 0.00443f
C1289 XA20.XA2a.MN0.D XA3.XA1.XA2.MP0.D 0.227f
C1290 XA20.XA2.MN1.D a_23600_44804# 0.0523f
C1291 XA1.XA4.MN0.G a_3440_42340# 7.97e-19
C1292 XA3.XA3.MN0.G a_9848_43396# 7.98e-19
C1293 XA2.XA1.XA5.MN2.D a_5960_44100# 0.126f
C1294 a_8480_45508# EN 3.34e-19
C1295 SARN XA5.XA6.MP0.G 0.0424f
C1296 XA8.XA7.MP0.G a_19928_51140# 0.0661f
C1297 a_8480_51140# a_9848_51140# 8.89e-19
C1298 AVDD a_4808_47268# 0.00125f
C1299 XA2.XA1.XA5.MN2.G D<7> 0.691f
C1300 XB2.XA4.MP0.D XDAC2.XC1.XRES16.B 0.0646f
C1301 XA3.XA3.MN0.G a_8480_40932# 0.00366f
C1302 EN XA1.XA1.XA4.MP1.D 0.0386f
C1303 XA0.XA1.XA5.MP0.D a_920_43396# 0.049f
C1304 AVDD a_18560_44100# 0.00125f
C1305 a_920_50436# VREF 0.0035f
C1306 XA4.XA6.MP0.D a_11000_50084# 0.049f
C1307 XA3.XA1.XA5.MN2.G a_7328_48324# 7.1e-20
C1308 XA4.XA1.XA5.MN2.G a_5960_48324# 7.1e-20
C1309 D<8> li_14804_25524# 3.5e-20
C1310 XA3.XA1.XA4.MN0.D a_7328_42340# 2.16e-19
C1311 XA3.XA1.XA4.MP0.D a_8480_42340# 2.16e-19
C1312 EN a_920_40228# 0.0674f
C1313 a_13520_48676# a_14888_48676# 8.89e-19
C1314 XA4.XA1.XA5.MN2.G a_9848_45156# 1e-19
C1315 D<6> a_5960_45508# 0.00436f
C1316 XA3.XA4.MN0.D XA20.XA3a.MN0.D 0.0699f
C1317 AVDD a_4808_41636# 0.00125f
C1318 XA4.XA6.MP0.G XA2.XA3.MN0.G 0.594f
C1319 VREF a_2288_47620# 0.0671f
C1320 D<2> a_16040_45860# 0.0774f
C1321 XA1.XA6.MP0.G a_2288_46564# 5.5e-19
C1322 a_18560_54308# XA8.XA11.MN1.G 6.78e-19
C1323 AVDD XA1.XA11.MP0.D 0.176f
C1324 a_4808_53956# XA3.XA11.MN1.G 0.0224f
C1325 XA20.XA12.MP0.G a_19928_53604# 0.00224f
C1326 a_18560_41284# XA7.XA1.XA1.MN0.D 0.00224f
C1327 a_7328_41284# a_7328_40932# 0.0109f
C1328 VREF a_16040_44452# 0.0182f
C1329 XA5.XA6.MP0.G a_13520_43748# 7.76e-20
C1330 D<3> a_13520_43044# 6.49e-19
C1331 XA1.XA6.MP0.G XA1.XA1.XA2.MP0.D 0.0106f
C1332 XA5.XA4.MN0.G a_12368_45860# 2.12e-19
C1333 AVDD a_13808_1390# 0.00159f
C1334 a_8480_46916# a_9848_46916# 8.89e-19
C1335 D<7> XA1.XA1.XA4.MN1.D 0.00188f
C1336 XA6.XA1.XA5.MN2.G a_14888_42692# 0.0739f
C1337 XA2.XA11.MN1.G XA1.XA8.MP0.D 2.37e-19
C1338 a_7328_52900# a_7328_52548# 0.0109f
C1339 a_18560_52900# XA7.XA10.MP0.G 0.0665f
C1340 XA7.XA10.MP0.D a_18560_52548# 0.00316f
C1341 AVDD a_23600_51140# 0.00181f
C1342 CK_SAMPLE a_19928_51492# 0.00264f
C1343 a_9560_3150# XB1.XA1.MP0.D 0.00203f
C1344 SARN a_13808_686# 2.97e-20
C1345 XA5.XA1.XA5.MN2.G a_12368_39876# 0.00278f
C1346 D<7> a_2288_40228# 3.45e-20
C1347 XA6.XA3.MN0.G EN 0.00979f
C1348 XA20.XA3a.MN0.D a_920_43396# 0.00213f
C1349 AVDD XDAC2.XC1.XRES16.B 3.93e-19
C1350 XA3.XA1.XA5.MN2.D XA4.XA1.XA5.MN2.D 0.00869f
C1351 a_11000_45508# a_11000_45156# 0.0109f
C1352 D<3> a_12368_40580# 4.18e-20
C1353 XA3.XA6.MP0.G a_8480_41284# 3.97e-20
C1354 XA3.XA4.MN0.G a_8480_43044# 0.0409f
C1355 XA3.XA7.MP0.D a_8480_51140# 0.00388f
C1356 CK_SAMPLE a_13520_49028# 7.31e-19
C1357 AVDD a_3440_48324# 0.00131f
C1358 XA3.XA8.MP0.D a_8480_51492# 0.00224f
C1359 a_18560_51844# a_18560_51492# 0.0109f
C1360 li_9184_29004# li_9184_28392# 0.00271f
C1361 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES2.B 0.0307f
C1362 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES16.B 0.0381f
C1363 XDAC1.XC0.XRES1A.B XDAC1.XC64b<1>.XRES1A.B 0.00444f
C1364 XA2.XA6.MP0.G XDAC2.XC0.XRES16.B 2.19e-20
C1365 XA20.XA3a.MN0.D a_n232_40932# 0.0739f
C1366 XA20.XA2a.MN0.D a_7328_41988# 0.00302f
C1367 XA4.XA1.XA5.MP1.D a_9848_43748# 2.16e-19
C1368 XA4.XA1.XA5.MN1.D a_11000_43748# 2.16e-19
C1369 XA0.XA6.MP2.G li_9184_20208# 3.5e-20
C1370 EN a_22448_43748# 5.7e-20
C1371 a_23600_44100# a_23600_43748# 0.0109f
C1372 AVDD a_7328_45156# 0.356f
C1373 a_23600_51140# XA20.XA3.MN0.D 3.51e-20
C1374 XA4.XA1.XA5.MN2.G XA3.XA4.MN0.D 0.198f
C1375 XA7.XA1.XA5.MN2.G VREF 0.704f
C1376 D<0> XA8.XA6.MN0.D 0.00148f
C1377 XDAC2.XC32a<0>.XRES16.B li_14804_13248# 0.00117f
C1378 XA1.XA4.MN0.D li_9184_9768# 0.00504f
C1379 XA0.XA4.MN0.D XDAC1.XC64a<0>.XRES1A.B 2.23e-21
C1380 a_n232_42692# a_920_42692# 0.00133f
C1381 D<2> a_14888_46916# 0.00249f
C1382 D<5> XA1.XA3.MN0.G 0.0259f
C1383 a_7328_49380# a_7328_49028# 0.0109f
C1384 XA0.XA6.MP2.G a_920_46564# 0.0695f
C1385 XA4.XA1.XA5.MN2.G a_7328_46212# 0.00363f
C1386 AVDD a_14888_42692# 0.00125f
C1387 VREF a_920_48676# 0.0191f
C1388 XA7.XA4.MN0.D a_17408_49028# 0.154f
C1389 AVDD a_13520_54308# 0.00166f
C1390 SARP XDAC1.X16ab.XRES8.B 27.7f
C1391 VREF a_16040_45508# 0.0556f
C1392 XA7.XA6.MP0.G a_17408_44804# 5.5e-19
C1393 XA2.XA1.XA5.MN2.G a_3440_43396# 2.66e-19
C1394 XA0.XA7.MP0.G a_4808_43396# 7.1e-20
C1395 XA8.XA1.XA5.MN2.G XA8.XA1.XA2.MP0.D 0.126f
C1396 XA0.XA6.MP2.G XA0.XA1.XA5.MP0.D 7.42e-19
C1397 a_2288_47620# a_2288_47268# 0.0109f
C1398 AVDD a_11000_39876# 0.44f
C1399 XA5.XA6.MP0.G SARP 0.0253f
C1400 a_18560_53252# a_19928_53252# 8.89e-19
C1401 AVDD a_5960_51844# 0.387f
C1402 XA0.XA12.MP0.D XA0.XA9.MN1.G 0.00116f
C1403 XA6.XA11.MN1.G a_12368_52548# 7.25e-20
C1404 a_21080_40228# a_22448_40228# 8.89e-19
C1405 D<2> XA6.XA1.XA1.MN0.S 0.018f
C1406 a_22448_46212# a_22448_45860# 0.0109f
C1407 XA8.XA4.MN0.G XA8.XA1.XA5.MN1.D 0.0242f
C1408 XA2.XA4.MN0.G a_4808_43748# 0.0157f
C1409 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MP1.D 0.148f
C1410 XA7.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.D 0.0326f
C1411 XA0.XA7.MP0.G a_3440_40932# 0.00631f
C1412 XA2.XA1.XA5.MN2.G a_2288_40932# 0.0245f
C1413 XA5.XA9.MN1.G XA5.XA8.MP0.D 0.0132f
C1414 a_22448_55364# VREF 0.0015f
C1415 XA20.XA4.MN0.D XA8.XA7.MP0.G 8.03e-19
C1416 a_5960_52548# XA3.XA1.XA5.MN2.G 1.75e-19
C1417 a_21080_52196# XA8.XA7.MP0.D 0.0658f
C1418 XA2.XA7.MP0.D XA3.XA7.MP0.D 0.00435f
C1419 AVDD XA1.XA4.MN0.D 2.65f
C1420 CK_SAMPLE a_13520_50084# 0.167f
C1421 XA2.XA9.MN1.G a_3440_51492# 2.84e-19
C1422 a_9848_52196# a_9848_51844# 0.0109f
C1423 a_11000_n18# a_12368_n18# 8.89e-19
C1424 XA2.XA4.MN0.D a_5960_40228# 9.14e-20
C1425 D<7> XDAC1.XC0.XRES16.B 5.78e-20
C1426 a_7328_44452# EN 0.00173f
C1427 a_16040_44452# a_16040_44100# 0.0109f
C1428 XA20.XA2a.MN0.D XA6.XA1.XA4.MN1.D 0.0128f
C1429 XA3.XA6.MN2.D a_8480_50788# 0.0488f
C1430 XA2.XA1.XA5.MN2.G XA2.XA6.MP0.G 0.00254f
C1431 AVDD a_4808_46212# 0.00125f
C1432 a_23600_51140# a_23600_50788# 0.0109f
C1433 XA20.XA2a.MN0.D a_13520_40228# 2.1e-19
C1434 XA3.XA1.XA2.MP0.D a_7328_42692# 7.68e-20
C1435 a_16040_43396# a_16040_43044# 0.0109f
C1436 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES16.B 0.0269f
C1437 XA4.XA1.XA5.MN2.G a_5960_47268# 7.1e-20
C1438 XA3.XA1.XA5.MN2.G a_7328_47268# 7.1e-20
C1439 AVDD XA8.XA1.XA5.MP0.D 0.143f
C1440 a_12368_49732# a_13520_49732# 0.00133f
C1441 a_920_49732# XA0.XA4.MN0.D 0.0658f
C1442 XA0.XA6.MP2.G XA20.XA3a.MN0.D 0.0701f
C1443 D<4> a_9848_47972# 5.43e-19
C1444 a_2288_42340# XA1.XA1.XA1.MN0.S 1.34e-19
C1445 a_2288_41988# a_2288_41636# 0.0109f
C1446 D<2> a_16040_44804# 2.36e-19
C1447 a_14888_48324# a_14888_47972# 0.0109f
C1448 XA1.XA4.MN0.G a_3440_47972# 0.153f
C1449 XA6.XA4.MN0.G XA7.XA4.MN0.G 0.00869f
C1450 D<6> a_4808_44452# 5.24e-19
C1451 XA1.XA4.MN0.D a_2288_46564# 2.2e-19
C1452 VREF a_3440_46564# 7.39e-19
C1453 AVDD XA8.XA1.XA1.MN0.D 0.0421f
C1454 XA6.XA4.MN0.D XA6.XA3.MN0.G 0.00642f
C1455 XA7.XA1.XA5.MN2.G a_16040_44100# 0.00556f
C1456 a_n232_53604# XA0.XA11.MN1.G 0.0709f
C1457 XA7.XA11.MN1.G XA6.XA11.MP0.D 0.00856f
C1458 AVDD a_2288_52548# 0.405f
C1459 XA2.XA12.MP0.G a_4808_53252# 0.0661f
C1460 XA3.XA11.MN1.G a_5960_53252# 0.00648f
C1461 XA5.XA1.XA1.MN0.D a_13520_40228# 0.00155f
C1462 a_14888_40932# a_14888_40580# 0.0109f
C1463 VREF XA1.XA1.XA5.MP0.D 0.00202f
C1464 XA1.XA4.MN0.D XA1.XA1.XA2.MP0.D 0.0111f
C1465 XA3.XA1.XA5.MN2.G a_7328_41636# 4.13e-19
C1466 a_16040_46564# a_17408_46564# 8.89e-19
C1467 a_3440_46564# a_3440_46212# 0.0109f
C1468 XA5.XA4.MN0.G a_12368_44804# 5.54e-19
C1469 XA5.XA3.MN0.G a_12368_46212# 0.155f
C1470 XA20.XA10.MN1.D a_23600_51140# 0.00455f
C1471 CK_SAMPLE a_12368_50788# 0.00142f
C1472 a_19928_52548# XA8.XA9.MN1.G 0.0727f
C1473 AVDD XA0.XA6.MP0.D 0.144f
C1474 XB1.M1.G a_11000_1038# 0.163f
C1475 SAR_IP CK_SAMPLE_BSSW 0.0123f
C1476 XB1.XA0.MP0.D XB1.XA3.MN0.S 0.572f
C1477 XB2.XA0.MP0.D a_14960_1742# 0.135f
C1478 a_13808_2094# XB2.XA3.MN0.S 3.29e-19
C1479 SAR_IN a_13808_686# 5.55e-19
C1480 XB2.M1.G a_14960_1390# 5.05e-19
C1481 XA20.XA3a.MN0.D a_16040_42692# 0.00443f
C1482 a_9848_44804# a_11000_44804# 0.00133f
C1483 a_23600_45156# a_23600_44804# 0.0109f
C1484 XA6.XA6.MP0.G a_12368_40580# 3.3e-20
C1485 XA1.XA4.MN0.G a_2288_42340# 1.28e-19
C1486 XA7.XA4.MN0.G XA7.XA1.XA4.MN0.D 0.00331f
C1487 XA3.XA3.MN0.G a_8480_43396# 0.00348f
C1488 XA2.XA1.XA5.MN2.D a_4808_44100# 0.0877f
C1489 a_7328_45508# EN 1.42e-19
C1490 SARN li_14804_25524# 0.00103f
C1491 AVDD a_3440_47268# 0.00125f
C1492 XA0.XA7.MP0.G D<7> 0.0713f
C1493 XA6.XA9.MN1.G XA6.XA6.MP0.D 0.0618f
C1494 a_12368_52900# VREF 0.00396f
C1495 XB1.XA4.MP0.D XDAC1.XC1.XRES1A.B 0.379f
C1496 XDAC2.X16ab.XRES16.B XDAC2.X16ab.XRES1A.B 0.454f
C1497 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES1A.B 0.00405f
C1498 EN XA0.XA1.XA4.MP1.D 0.0393f
C1499 XA20.XA2a.MN0.D a_22448_41284# 0.00107f
C1500 XA0.XA1.XA5.MP0.D a_n232_43396# 2.16e-19
C1501 XA0.XA1.XA5.MN0.D a_920_43396# 2.16e-19
C1502 a_13520_43748# a_13520_43396# 0.0109f
C1503 AVDD a_17408_44100# 0.359f
C1504 XA0.XA6.MP0.G a_920_49732# 0.101f
C1505 XA0.XA6.MN0.D a_n232_49732# 0.00176f
C1506 XA3.XA1.XA5.MN2.G a_5960_48324# 0.00455f
C1507 XDAC2.XC64a<0>.XRES16.B XDAC2.XC1.XRES16.B 0.0114f
C1508 li_14804_8736# li_14804_8124# 0.00271f
C1509 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES8.B 0.0228f
C1510 XA3.XA3.MN0.G li_14804_26136# 0.00504f
C1511 SARP a_9560_3854# 0.00146f
C1512 XA0.XA1.XA2.MP0.D a_920_40932# 4.25e-20
C1513 XA3.XA1.XA4.MP0.D a_7328_42340# 0.049f
C1514 a_19928_42692# a_19928_42340# 0.0109f
C1515 EN a_n232_40228# 0.0708f
C1516 D<6> a_4808_45508# 0.0031f
C1517 XA7.XA4.MN0.D a_18560_47972# 0.0788f
C1518 XA2.XA4.MN0.D XA20.XA3a.MN0.D 0.0705f
C1519 a_920_48676# a_920_48324# 0.0109f
C1520 XA4.XA1.XA5.MN2.G a_8480_45156# 1.95e-19
C1521 AVDD a_3440_41636# 0.00125f
C1522 XA4.XA6.MP0.G XA1.XA3.MN0.G 0.027f
C1523 VREF a_920_47620# 0.0671f
C1524 D<2> a_14888_45860# 0.0675f
C1525 a_17408_54308# XA8.XA11.MN1.G 8.3e-19
C1526 a_16040_53956# a_17408_53956# 8.89e-19
C1527 AVDD XA0.XA11.MP0.D 0.19f
C1528 XA2.XA1.XA1.MN0.S a_5960_40580# 0.0318f
C1529 XA7.XA1.XA1.MP2.D a_17408_40932# 0.00176f
C1530 SARP li_9184_15084# 0.00103f
C1531 XA5.XA6.MP0.G a_12368_43748# 5.5e-19
C1532 VREF a_14888_44452# 7.12e-19
C1533 D<3> a_12368_43044# 7.77e-20
C1534 a_21080_47268# a_21080_46916# 0.0109f
C1535 D<7> XA1.XA1.XA4.MP1.D 7.43e-19
C1536 XA6.XA1.XA5.MN2.G a_13520_42692# 1.95e-19
C1537 a_13520_53252# XA5.XA9.MN1.G 5.25e-19
C1538 a_17408_52900# XA7.XA10.MP0.G 0.0674f
C1539 XA0.XA10.MP0.G XA1.XA10.MP0.G 0.00217f
C1540 XA7.XA10.MP0.D a_17408_52548# 0.00224f
C1541 AVDD a_22448_51140# 0.569f
C1542 CK_SAMPLE a_18560_51492# 6.45e-19
C1543 a_13808_3150# a_14960_3150# 0.00133f
C1544 XB1.XA2.MN0.G XB1.XA1.MN0.D 0.0103f
C1545 a_8408_3150# XB1.XA1.MP0.D 4.43e-19
C1546 XA8.XA3.MN0.G a_21080_44100# 0.00245f
C1547 XA1.XA3.MN0.G XA1.XA1.XA5.MN1.D 0.00103f
C1548 XA5.XA3.MN0.G EN 0.00979f
C1549 SARN a_12368_686# 0.0353f
C1550 XA7.XA6.MP0.G XA6.XA1.XA1.MN0.S 0.0022f
C1551 XA5.XA1.XA5.MN2.G a_11000_39876# 0.00285f
C1552 XA20.XA3a.MN0.D a_n232_43396# 0.0736f
C1553 AVDD XDAC1.XC1.XRES16.B 5.34e-19
C1554 XA3.XA6.MP0.G a_7328_41284# 4.24e-19
C1555 XA3.XA4.MN0.G a_7328_43044# 0.0222f
C1556 a_7328_51844# XA4.XA1.XA5.MN2.G 8.87e-19
C1557 XA0.XA9.MN1.G a_920_50788# 0.00281f
C1558 XA3.XA7.MP0.D a_7328_51140# 0.00224f
C1559 CK_SAMPLE a_12368_49028# 3.27e-19
C1560 XA3.XA8.MP0.D a_7328_51492# 0.00224f
C1561 a_n232_51492# a_920_51492# 0.00133f
C1562 AVDD a_2288_48324# 0.359f
C1563 XA20.XA2a.MN0.D a_5960_41988# 0.00302f
C1564 XA1.XA1.XA5.MN2.D a_2288_42692# 7.44e-20
C1565 XA20.XA3a.MN0.D XA8.XA1.XA1.MP1.D 0.0093f
C1566 XA4.XA1.XA5.MN1.D a_9848_43748# 0.0494f
C1567 EN a_21080_43748# 0.166f
C1568 a_12368_50436# a_13520_50436# 0.00133f
C1569 a_920_50436# XA0.XA6.MP0.G 0.0662f
C1570 AVDD a_5960_45156# 0.356f
C1571 XA8.XA7.MP0.G a_22448_49732# 0.00104f
C1572 a_11000_50788# XA4.XA6.MP0.G 1.34e-19
C1573 XA3.XA1.XA5.MN2.G XA3.XA4.MN0.D 0.069f
C1574 XA4.XA1.XA5.MN2.G XA2.XA4.MN0.D 6.95e-19
C1575 XA6.XA1.XA5.MN2.G VREF 0.704f
C1576 D<0> XA8.XA6.MP0.G 0.421f
C1577 a_n232_50436# XA0.XA6.MN0.D 0.00176f
C1578 XA1.XA1.XA2.MP0.D a_3440_41636# 0.00316f
C1579 XA5.XA1.XA2.MP0.D a_13520_41988# 0.0568f
C1580 XA4.XA1.XA4.MP1.D a_11000_42692# 0.049f
C1581 a_23600_43044# a_23600_42692# 0.0109f
C1582 D<5> D<8> 0.0323f
C1583 XA8.XA6.MP0.G XA8.XA4.MN0.G 0.0052f
C1584 XA1.XA6.MP0.G XA20.XA3a.MN0.D 0.0676f
C1585 a_18560_49380# a_19928_49380# 8.89e-19
C1586 XA0.XA6.MP2.G a_n232_46564# 0.0551f
C1587 XA3.XA1.XA5.MN2.G a_7328_46212# 7.1e-20
C1588 XA4.XA1.XA5.MN2.G a_5960_46212# 7.1e-20
C1589 D<6> XA3.XA3.MN0.G 0.144f
C1590 AVDD a_13520_42692# 0.00125f
C1591 XA0.XA4.MN0.D a_920_48676# 0.154f
C1592 VREF a_n232_48676# 1.3e-19
C1593 AVDD a_12368_54308# 0.448f
C1594 XA20.XA1.MN0.D a_23600_40932# 0.0562f
C1595 XA3.XA1.XA1.MN0.S XA4.XA1.XA1.MN0.S 0.00217f
C1596 a_21080_41636# XA8.XA1.XA1.MP2.D 0.00176f
C1597 a_9848_41636# a_9848_41284# 0.0109f
C1598 XA4.XA4.MN0.G a_11000_46916# 0.0678f
C1599 XA2.XA1.XA5.MN2.G a_2288_43396# 0.00442f
C1600 XA0.XA7.MP0.G a_3440_43396# 0.00518f
C1601 D<4> a_11000_43748# 7.76e-20
C1602 XA8.XA1.XA5.MN2.G XA7.XA1.XA5.MN0.D 7.2e-19
C1603 XA7.XA1.XA5.MN2.G XA8.XA1.XA2.MP0.D 1.74e-19
C1604 XA0.XA6.MP2.G XA0.XA1.XA5.MN0.D 0.00188f
C1605 a_13520_47620# a_14888_47620# 8.89e-19
C1606 AVDD a_9848_39876# 0.00131f
C1607 XA3.XA11.MP0.D a_7328_52900# 0.00176f
C1608 a_8480_53252# XA3.XA10.MP0.D 0.0676f
C1609 a_n232_53252# a_n232_52900# 0.0109f
C1610 AVDD a_4808_51844# 0.00166f
C1611 XA5.XA11.MN1.G a_13520_52548# 0.00103f
C1612 a_8480_40228# a_8480_39876# 0.0109f
C1613 a_8480_45860# a_9848_45860# 8.89e-19
C1614 XA5.XA3.MN0.G a_13520_45156# 0.0805f
C1615 XA20.XA3a.MN0.D a_18560_44100# 5.04e-20
C1616 D<6> a_5960_41284# 7.76e-20
C1617 XA7.XA1.XA5.MN2.G XA7.XA1.XA1.MP1.D 6.68e-19
C1618 XA0.XA7.MP0.G a_2288_40932# 0.0013f
C1619 XA2.XA4.MN0.D XA2.XA1.XA4.MP1.D 9.69e-19
C1620 XA1.XA9.MN1.G a_4808_51492# 2.84e-19
C1621 a_19928_52196# XA8.XA7.MP0.D 0.0678f
C1622 AVDD VREF 69.8f
C1623 CK_SAMPLE a_12368_50084# 0.00848f
C1624 a_14960_334# a_14960_n18# 0.0109f
C1625 XA2.XA4.MN0.D a_4808_40228# 9.25e-20
C1626 XA0.XA6.MP2.G li_9184_30648# 0.00508f
C1627 a_5960_44452# EN 0.00173f
C1628 a_2288_44100# a_3440_44100# 0.00133f
C1629 XA20.XA3a.MN0.D a_4808_41636# 0.00547f
C1630 SARN XDAC2.XC32a<0>.XRES4.B 13.9f
C1631 XA20.XA2a.MN0.D XA5.XA1.XA4.MN1.D 0.0128f
C1632 D<1> XA7.XA6.MN2.D 1.59e-19
C1633 XA8.XA7.MP0.G a_22448_50436# 0.00126f
C1634 XA5.XA9.MN1.G a_13520_49380# 4.23e-20
C1635 AVDD a_3440_46212# 0.00125f
C1636 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES8.B 0.471f
C1637 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES2.B 0.0136f
C1638 a_2288_43044# a_3440_43044# 0.00133f
C1639 XA0.XA6.MP0.G li_14804_9768# 1.85e-20
C1640 XA0.XA4.MN0.D XDAC1.XC128b<2>.XRES1A.B 0.00405f
C1641 EN a_17408_42340# 0.159f
C1642 D<1> XA7.XA4.MN0.G 0.26f
C1643 XA3.XA1.XA5.MN2.G a_5960_47268# 0.00363f
C1644 AVDD XA8.XA1.XA5.MN0.D 0.00912f
C1645 XA4.XA6.MP0.G a_11000_49028# 0.0307f
C1646 XA0.XA6.MP0.G a_920_48676# 0.0881f
C1647 XA8.XA6.MP0.G a_21080_49380# 0.0781f
C1648 a_n232_49732# XA0.XA4.MN0.D 0.0675f
C1649 XA20.XA3.MN0.D VREF 6.24e-19
C1650 a_13520_41988# a_14888_41988# 8.89e-19
C1651 XA1.XA4.MN0.G a_2288_47972# 0.155f
C1652 VREF a_2288_46564# 0.0175f
C1653 AVDD XA7.XA1.XA1.MN0.D 0.0357f
C1654 XA7.XA1.XA5.MN2.G a_14888_44100# 2.31e-19
C1655 D<2> a_14888_44804# 5.24e-19
C1656 a_11000_53604# a_12368_53604# 8.89e-19
C1657 AVDD a_920_52548# 0.405f
C1658 CK_SAMPLE XA20.XA9.MP0.D 0.0123f
C1659 XA3.XA11.MN1.G a_4808_53252# 2.82e-19
C1660 a_920_40580# a_2288_40580# 8.89e-19
C1661 XA0.XA11.MN1.G XB2.XA4.MP0.D 7.2e-20
C1662 XA3.XA1.XA5.MN2.G a_5960_41636# 0.0756f
C1663 XA1.XA10.MP0.G XA1.XA7.MP0.D 0.0601f
C1664 XA7.XA10.MP0.G a_18560_52196# 0.0131f
C1665 CK_SAMPLE a_11000_50788# 0.00142f
C1666 a_7328_52548# a_7328_52196# 0.0109f
C1667 AVDD XA0.XA6.MN0.D 3.13e-19
C1668 XA20.XA10.MN1.D a_22448_51140# 1.97e-19
C1669 a_9560_1742# a_11000_1742# 8e-19
C1670 XB1.XA4.MP0.D a_8408_1038# 0.00161f
C1671 XB1.M1.G a_9560_1038# 0.00112f
C1672 XB2.XA0.MP0.D a_13808_1742# 0.0781f
C1673 SAR_IN a_12368_686# 0.0598f
C1674 XB2.M1.G a_13808_1390# 0.0015f
C1675 XA20.XA3a.MN0.D a_14888_42692# 0.0099f
C1676 XA8.XA1.XA5.MN2.D a_21080_44452# 0.158f
C1677 a_5960_45508# EN 1.42e-19
C1678 XA6.XA9.MN1.G XA6.XA6.MN0.D 0.0615f
C1679 a_7328_51140# a_8480_51140# 0.00133f
C1680 XA8.XA1.XA5.MN2.G a_18560_51140# 0.0677f
C1681 AVDD a_2288_47268# 0.356f
C1682 XA0.XA7.MP0.G XA0.XA6.MP2.D 0.00313f
C1683 a_11000_52900# VREF 0.00396f
C1684 XA0.XA9.MN1.G a_920_50084# 0.00281f
C1685 XA4.XA7.MP0.D a_9848_50436# 1.37e-19
C1686 EN XA0.XA1.XA4.MN1.D 0.0134f
C1687 XA1.XA6.MP0.G XDAC2.XC128b<2>.XRES16.B 4.21e-20
C1688 XA20.XA2a.MN0.D a_21080_41284# 0.0672f
C1689 XA0.XA1.XA5.MN0.D a_n232_43396# 0.0474f
C1690 XA4.XA6.MN0.D a_9848_50084# 0.0488f
C1691 XA4.XA6.MP0.G a_11000_50084# 0.159f
C1692 AVDD a_16040_44100# 0.359f
C1693 XA0.XA6.MP0.G a_n232_49732# 0.00239f
C1694 XA8.XA7.MP0.G a_22448_48676# 8.22e-19
C1695 XA8.XA6.MP0.G XA20.XA3a.MN0.G 0.00435f
C1696 a_5960_43044# XA2.XA1.XA1.MN0.S 4.06e-20
C1697 SARP a_8408_3854# 2.37e-19
C1698 D<8> XDAC2.X16ab.XRES4.B 4.06e-21
C1699 XA3.XA1.XA5.MN2.G a_8480_45156# 1e-19
C1700 XA4.XA1.XA5.MN2.G a_7328_45156# 0.00486f
C1701 VREF a_n232_47620# 7.12e-19
C1702 XA7.XA4.MN0.D a_17408_47972# 0.0546f
C1703 XA1.XA4.MN0.D XA20.XA3a.MN0.D 0.0699f
C1704 a_12368_48676# a_13520_48676# 0.00133f
C1705 XA3.XA6.MP0.G XA3.XA3.MN0.G 3.29f
C1706 AVDD a_2288_41636# 0.404f
C1707 XA4.XA6.MP0.G D<8> 0.0334f
C1708 XA0.XA4.MN0.D a_920_47620# 0.00498f
C1709 D<2> a_13520_45860# 1.06e-19
C1710 AVDD XA0.XA11.MN1.G 9.55f
C1711 a_3440_53956# XA1.XA12.MP0.G 0.0688f
C1712 a_4808_53956# XA2.XA11.MN1.G 7.59e-19
C1713 a_18560_54308# XA7.XA11.MN1.G 0.00123f
C1714 XA2.XA1.XA1.MN0.S a_4808_40580# 0.00155f
C1715 XA7.XA1.XA1.MN0.S a_17408_40932# 0.0271f
C1716 a_17408_41284# XA7.XA1.XA1.MP1.D 0.00176f
C1717 a_5960_41284# a_5960_40932# 0.0109f
C1718 XA4.XA4.MN0.G a_11000_45860# 2.12e-19
C1719 a_7328_46916# a_8480_46916# 0.00133f
C1720 XA6.XA1.XA5.MN2.G a_12368_42692# 0.00442f
C1721 XA5.XA1.XA5.MN2.G a_13520_42692# 0.0755f
C1722 VREF a_13520_44452# 7.12e-19
C1723 XA6.XA11.MN1.G a_13520_51844# 1.13e-19
C1724 XA0.XA10.MP0.D XA0.XA9.MN1.G 0.00406f
C1725 a_5960_52900# a_5960_52548# 0.0109f
C1726 AVDD a_21080_51140# 0.382f
C1727 CK_SAMPLE a_17408_51492# 5.02e-19
C1728 XA0.XA12.MP0.D XA1.XA8.MP0.D 6.42e-19
C1729 XB1.XA2.MN0.G XB1.XA1.MP0.D 0.00383f
C1730 XB2.XA2.MN0.G a_14960_3150# 0.0731f
C1731 XA8.XA3.MN0.G a_19928_44100# 0.00441f
C1732 XA4.XA3.MN0.G EN 0.00979f
C1733 XA0.XA4.MN0.D a_920_41988# 9.14e-20
C1734 SARN a_11000_686# 5.3e-20
C1735 XA20.XA3a.MN0.D XA8.XA1.XA5.MP0.D 0.0273f
C1736 XA2.XA1.XA5.MN2.D XA3.XA1.XA5.MN2.D 0.00869f
C1737 a_21080_45508# XA8.XA1.XA5.MN2.D 0.0659f
C1738 a_9848_45508# a_9848_45156# 0.0109f
C1739 XA0.XA9.MN1.G a_n232_50788# 0.015f
C1740 XA20.XA10.MN1.D VREF 0.00546f
C1741 a_17408_51844# a_17408_51492# 0.0109f
C1742 XA5.XA9.MN1.G XA5.XA6.MN2.D 0.126f
C1743 SARN D<5> 0.027f
C1744 AVDD a_920_48324# 0.359f
C1745 CK_SAMPLE a_11000_49028# 3.27e-19
C1746 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES8.B 0.471f
C1747 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES2.B 0.0136f
C1748 XA8.XA1.XA5.MN1.D XA8.XA1.XA5.MP1.D 0.00918f
C1749 XA20.XA2a.MN0.D a_4808_41988# 0.0844f
C1750 XA20.XA3a.MN0.D XA8.XA1.XA1.MN0.D 0.0616f
C1751 XA0.XA6.MP2.G XDAC1.XC128b<2>.XRES16.B 3.84e-19
C1752 a_18560_44452# XA7.XA1.XA2.MP0.D 5.16e-20
C1753 a_8480_44100# XA3.XA1.XA2.MP0.D 2.92e-19
C1754 EN a_19928_43748# 0.00532f
C1755 a_22448_44100# a_22448_43748# 0.0109f
C1756 AVDD a_4808_45156# 0.00125f
C1757 XA8.XA7.MP0.G a_21080_49732# 0.00457f
C1758 a_9848_50788# XA4.XA6.MP0.G 1.75e-20
C1759 XA3.XA1.XA5.MN2.G XA2.XA4.MN0.D 0.123f
C1760 XA5.XA1.XA5.MN2.G VREF 0.704f
C1761 a_n232_50436# XA0.XA6.MP0.G 3.02e-20
C1762 XDAC2.XC32a<0>.XRES4.B XDAC2.XC64a<0>.XRES4.B 0.00284f
C1763 li_14804_13860# li_14804_13248# 0.00271f
C1764 XDAC1.XC32a<0>.XRES16.B li_9184_13248# 0.00117f
C1765 EN a_7328_41284# 0.00564f
C1766 XA0.XA4.MN0.D li_9184_9768# 1.85e-20
C1767 XA1.XA4.MN0.D XDAC1.XC64a<0>.XRES16.B 0.0269f
C1768 XA4.XA1.XA4.MP1.D a_9848_42692# 2.16e-19
C1769 XA4.XA1.XA4.MN1.D a_11000_42692# 2.16e-19
C1770 XA1.XA1.XA2.MP0.D a_2288_41636# 0.00224f
C1771 XA5.XA1.XA2.MP0.D a_12368_41988# 0.0219f
C1772 XA0.XA6.MP0.G a_920_47620# 6.35e-19
C1773 a_5960_49380# a_5960_49028# 0.0109f
C1774 XA8.XA7.MP0.G XA20.XA2a.MN0.D 0.285f
C1775 XA3.XA1.XA5.MN2.G a_5960_46212# 0.00363f
C1776 D<6> XA2.XA3.MN0.G 1.02f
C1777 AVDD a_12368_42692# 0.358f
C1778 XA0.XA4.MN0.D a_n232_48676# 0.158f
C1779 XA6.XA4.MN0.D a_16040_49028# 0.154f
C1780 DONE XA20.XA11.MP0.D 0.0128f
C1781 AVDD a_11000_54308# 0.447f
C1782 SARP li_9184_25524# 0.00103f
C1783 a_21080_41636# XA8.XA1.XA1.MN0.S 0.0694f
C1784 XA3.XA1.XA1.MN0.S XA3.XA1.XA1.MP2.D 0.0708f
C1785 XA20.XA1.MN0.D a_22448_40932# 3.45e-19
C1786 XA8.XA1.XA5.MN2.G XA7.XA1.XA5.MP0.D 0.00353f
C1787 XA0.XA6.MP2.G XA0.XA1.XA2.MP0.D 0.0131f
C1788 a_920_47620# a_920_47268# 0.0109f
C1789 XA4.XA4.MN0.G a_9848_46916# 0.0869f
C1790 D<4> a_9848_43748# 6.49e-19
C1791 AVDD a_8480_39876# 0.00131f
C1792 a_17408_53252# a_18560_53252# 0.00133f
C1793 a_7328_53252# XA3.XA10.MP0.D 0.0677f
C1794 AVDD a_3440_51844# 0.00166f
C1795 XA5.XA11.MN1.G a_12368_52548# 0.00135f
C1796 a_19928_40228# a_21080_40228# 0.00133f
C1797 SARN a_23600_39876# 9.45e-19
C1798 a_21080_46212# a_21080_45860# 0.0109f
C1799 XA7.XA4.MN0.G XA7.XA1.XA5.MN1.D 0.0242f
C1800 XA1.XA4.MN0.G a_3440_43748# 0.0157f
C1801 XA5.XA3.MN0.G a_12368_45156# 0.0546f
C1802 D<6> a_4808_41284# 6.49e-19
C1803 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MP1.D 0.144f
C1804 XA0.XA7.MP0.G a_920_40932# 0.0256f
C1805 XA4.XA6.MP0.G a_11000_42340# 5.5e-19
C1806 XA2.XA4.MN0.D XA2.XA1.XA4.MN1.D 9.9e-19
C1807 XA0.XA6.MP0.G a_920_41988# 5.5e-19
C1808 XA1.XA9.MN1.G a_3440_51492# 0.0118f
C1809 XA1.XA7.MP0.D XA2.XA7.MP0.D 0.00435f
C1810 AVDD XA0.XA4.MN0.D 2.65f
C1811 CK_SAMPLE a_11000_50084# 0.00848f
C1812 a_8480_52196# a_8480_51844# 0.0109f
C1813 XA8.XA9.MN0.D a_19928_51844# 0.00176f
C1814 XA8.XA9.MN1.G a_21080_51844# 6.57e-19
C1815 a_9560_n18# a_11000_n18# 8e-19
C1816 a_4808_44452# EN 0.00154f
C1817 a_14888_44452# a_14888_44100# 0.0109f
C1818 XA20.XA3a.MN0.D a_3440_41636# 0.00547f
C1819 XA20.XA2a.MN0.D XA5.XA1.XA4.MP1.D 0.0128f
C1820 XA4.XA1.XA5.MN2.D XA4.XA1.XA2.MP0.D 4.72e-19
C1821 XA4.XA4.MN0.G XA4.XA1.XA1.MN0.S 5.22e-20
C1822 XA3.XA6.MP2.D a_7328_50788# 0.049f
C1823 XA8.XA7.MP0.G a_21080_50436# 0.0046f
C1824 a_12368_51492# XA5.XA6.MP0.G 4.06e-20
C1825 XA5.XA9.MN1.G a_12368_49380# 2.54e-19
C1826 a_12368_52196# VREF 0.00396f
C1827 AVDD a_2288_46212# 0.356f
C1828 a_22448_51140# a_22448_50788# 0.0109f
C1829 D<1> XA7.XA6.MP2.D 0.0399f
C1830 a_14888_43396# a_14888_43044# 0.0109f
C1831 XA6.XA1.XA2.MP0.D XA6.XA1.XA4.MP1.D 4.34e-19
C1832 XA1.XA6.MP0.G li_14804_10380# 0.00504f
C1833 EN a_16040_42340# 0.159f
C1834 XA8.XA7.MP0.G a_22448_47620# 6.64e-19
C1835 AVDD XA8.XA1.XA2.MP0.D 0.27f
C1836 XA4.XA6.MP0.G a_9848_49028# 0.0137f
C1837 XA0.XA6.MP0.G a_n232_48676# 0.0651f
C1838 XA8.XA6.MP0.G a_19928_49380# 0.0547f
C1839 a_11000_49732# a_12368_49732# 8.89e-19
C1840 SARP a_11000_686# 0.0356f
C1841 a_920_41988# a_920_41636# 0.0109f
C1842 a_13520_48324# a_13520_47972# 0.0109f
C1843 XA5.XA4.MN0.G XA6.XA4.MN0.G 0.12f
C1844 VREF a_920_46564# 0.0175f
C1845 AVDD XA7.XA1.XA1.MP1.D 0.0599f
C1846 XA5.XA4.MN0.D XA5.XA3.MN0.G 0.00642f
C1847 D<5> SARP 0.0893f
C1848 XA6.XA1.XA5.MN2.G a_14888_44100# 0.0709f
C1849 XA2.XA11.MN1.G a_5960_53252# 0.0674f
C1850 XA5.XA12.MP0.G XA5.XA11.MP0.D 0.0612f
C1851 XA6.XA11.MN1.G XA6.XA11.MP0.D 0.0102f
C1852 AVDD a_n232_52548# 0.00166f
C1853 a_23600_54308# XA20.XA9.MP0.D 3.02e-20
C1854 CK_SAMPLE XA8.XA10.MP0.D 0.00163f
C1855 XA20.XA10.MN0.D a_23600_53604# 0.0465f
C1856 a_13520_40932# a_13520_40580# 0.0109f
C1857 XA3.XA1.XA5.MN2.G a_4808_41636# 0.128f
C1858 XA8.XA7.MP0.G a_22448_41988# 9.75e-19
C1859 VREF XA0.XA1.XA5.MP0.D 0.00202f
C1860 D<1> XA7.XA1.XA4.MN0.D 0.00144f
C1861 a_14888_46564# a_16040_46564# 0.00133f
C1862 a_2288_46564# a_2288_46212# 0.0109f
C1863 XA0.XA11.MN1.G XB2.XA4.MN0.D 7.05e-19
C1864 XA4.XA4.MN0.G a_11000_44804# 5.54e-19
C1865 XA4.XA3.MN0.G a_11000_46212# 0.155f
C1866 XA7.XA10.MP0.G a_17408_52196# 0.0441f
C1867 a_18560_52548# XA7.XA9.MN0.D 0.00176f
C1868 CK_SAMPLE a_9848_50788# 0.157f
C1869 AVDD XA0.XA6.MP0.G 5.93f
C1870 XA2.XA9.MN1.G XA3.XA9.MN1.G 0.00217f
C1871 XB1.M1.G a_8408_1038# 1.7e-19
C1872 a_14960_2094# a_14960_1742# 0.0109f
C1873 XB2.M1.G a_12368_1390# 0.0703f
C1874 XA20.XA3a.MN0.D a_13520_42692# 0.01f
C1875 XA5.XA6.MP0.G a_13520_40580# 7.76e-20
C1876 a_22448_45156# a_22448_44804# 0.0109f
C1877 a_8480_44804# a_9848_44804# 8.89e-19
C1878 XA20.XA2a.MN0.D XA2.XA1.XA2.MP0.D 0.223f
C1879 XA1.XA6.MP0.G a_3440_40228# 3.45e-20
C1880 XA0.XA4.MN0.G a_920_42340# 1.28e-19
C1881 XA1.XA1.XA5.MN2.D a_3440_44100# 0.0893f
C1882 XA8.XA1.XA5.MN2.D a_19928_44452# 0.153f
C1883 a_4808_45508# EN 3.34e-19
C1884 SARN XDAC2.X16ab.XRES4.B 13.9f
C1885 XA6.XA9.MN1.G XA6.XA6.MP0.G 0.0725f
C1886 XA8.XA1.XA5.MN2.G a_17408_51140# 0.0754f
C1887 AVDD a_920_47268# 0.356f
C1888 XA2.XA1.XA5.MN2.G XA0.XA6.MP2.G 3.47e-19
C1889 XA0.XA7.MP0.G XA0.XA6.MN2.D 6.33e-19
C1890 a_11000_51492# D<4> 2.41e-19
C1891 XA0.XA9.MN1.G a_n232_50084# 0.00969f
C1892 SARN XA4.XA6.MP0.G 0.0424f
C1893 XDAC1.X16ab.XRES16.B XDAC1.X16ab.XRES1A.B 0.454f
C1894 XDAC2.X16ab.XRES16.B li_14804_23688# 0.00117f
C1895 XA0.XA6.MP0.G li_14804_20208# 0.00504f
C1896 XA20.XA2a.MN0.D a_19928_41284# 0.0897f
C1897 XA4.XA1.XA5.MN0.D XA4.XA1.XA5.MP0.D 0.00918f
C1898 XA0.XA1.XA2.MP0.D a_n232_43396# 0.0945f
C1899 a_12368_43748# a_12368_43396# 0.0109f
C1900 a_22448_50788# VREF 0.0014f
C1901 D<5> a_8480_49028# 5.7e-19
C1902 XA4.XA6.MP0.G a_9848_50084# 6.4e-20
C1903 AVDD a_14888_44100# 0.00125f
C1904 XA8.XA7.MP0.G a_21080_48676# 0.00363f
C1905 D<1> a_18560_49380# 5.91e-19
C1906 XA8.XA6.MP0.G XA8.XA6.MP0.D 0.0392f
C1907 XDAC1.XC64a<0>.XRES16.B XDAC1.XC1.XRES16.B 0.0114f
C1908 li_9184_8736# li_9184_8124# 0.00271f
C1909 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES8.B 0.0228f
C1910 a_18560_42692# a_18560_42340# 0.0109f
C1911 XA2.XA1.XA4.MP0.D a_5960_42340# 0.049f
C1912 XA7.XA1.XA4.MP0.D XA7.XA1.XA4.MN0.D 0.00918f
C1913 SARP a_23600_39876# 0.00646f
C1914 XA3.XA3.MN0.G XDAC2.X16ab.XRES1B.B 0.00405f
C1915 EN a_22448_40580# 5.7e-20
C1916 XA4.XA1.XA5.MN2.G a_5960_45156# 7.1e-20
C1917 XA3.XA1.XA5.MN2.G a_7328_45156# 7.1e-20
C1918 VREF XA20.XA3a.MN0.D 0.13f
C1919 XA0.XA4.MN0.D a_n232_47620# 0.0396f
C1920 a_n232_48676# a_n232_48324# 0.0109f
C1921 XA6.XA6.MP0.G a_16040_46916# 5.5e-19
C1922 XA3.XA6.MP0.G XA2.XA3.MN0.G 0.0572f
C1923 AVDD a_920_41636# 0.404f
C1924 a_14888_53956# a_16040_53956# 0.00133f
C1925 AVDD a_23600_53604# 0.00154f
C1926 a_3440_53956# XA2.XA11.MN1.G 0.0225f
C1927 a_2288_53956# XA1.XA12.MP0.G 0.0674f
C1928 a_17408_54308# XA7.XA11.MN1.G 8.45e-19
C1929 SARP XDAC1.XC32a<0>.XRES4.B 13.9f
C1930 XA4.XA4.MN0.G a_9848_45860# 0.0146f
C1931 AVDD a_9560_1390# 0.00159f
C1932 a_9848_47268# XA4.XA3.MN0.G 2.69e-19
C1933 a_19928_47268# a_19928_46916# 0.0109f
C1934 XA5.XA1.XA5.MN2.G a_12368_42692# 1.97e-19
C1935 VREF a_12368_44452# 0.0182f
C1936 XA3.XA4.MN0.D a_8480_44452# 9.24e-20
C1937 a_16040_52900# XA6.XA10.MP0.G 0.0658f
C1938 XA6.XA10.MP0.D a_16040_52548# 0.00224f
C1939 AVDD a_19928_51140# 0.00166f
C1940 CK_SAMPLE a_16040_51492# 5.02e-19
C1941 a_9560_3502# XB1.XA1.MP0.D 2.12e-19
C1942 a_14960_3502# a_14960_3150# 0.0109f
C1943 XB2.XA2.MN0.G a_13808_3150# 0.0658f
C1944 XA4.XA1.XA5.MN2.G a_9848_39876# 0.00169f
C1945 XA3.XA3.MN0.G EN 0.0848f
C1946 XA0.XA4.MN0.D a_n232_41988# 9.25e-20
C1947 XA7.XA6.MP0.G XA5.XA1.XA1.MN0.S 5.61e-19
C1948 XA20.XA3a.MN0.D XA8.XA1.XA5.MN0.D 0.0353f
C1949 a_19928_45508# XA8.XA1.XA5.MN2.D 0.0674f
C1950 XA2.XA4.MN0.G a_5960_43044# 0.0222f
C1951 XA8.XA12.MP0.G VREF 0.0115f
C1952 XA2.XA8.MP0.D a_5960_51492# 0.00224f
C1953 a_5960_51844# XA3.XA1.XA5.MN2.G 8.87e-19
C1954 XA5.XA9.MN1.G XA5.XA6.MP2.D 0.0618f
C1955 AVDD a_n232_48324# 0.00131f
C1956 CK_SAMPLE a_9848_49028# 7.31e-19
C1957 XA8.XA7.MP0.D XA8.XA7.MP0.G 0.139f
C1958 XA2.XA7.MP0.D a_5960_51140# 0.00224f
C1959 XA20.XA3a.MN0.D XA7.XA1.XA1.MN0.D 0.0616f
C1960 XA3.XA1.XA5.MN1.D a_8480_43748# 0.0494f
C1961 XA20.XA2a.MN0.D a_3440_41988# 0.0861f
C1962 XA0.XA1.XA5.MN2.D a_920_42692# 7.44e-20
C1963 XA1.XA6.MP0.G XDAC2.XC0.XRES16.B 4.21e-20
C1964 EN a_18560_43748# 0.00532f
C1965 AVDD a_3440_45156# 0.00125f
C1966 a_11000_50436# a_12368_50436# 8.89e-19
C1967 XA4.XA1.XA5.MN2.G VREF 0.704f
C1968 XA2.XA1.XA5.MN2.G XA2.XA4.MN0.D 0.00344f
C1969 D<5> a_8480_50084# 5.7e-19
C1970 EN a_5960_41284# 0.00564f
C1971 XA4.XA1.XA4.MN1.D a_9848_42692# 0.0474f
C1972 a_22448_43044# a_22448_42692# 0.0109f
C1973 XA4.XA6.MP0.G a_11000_47972# 8.92e-19
C1974 a_17408_49380# a_18560_49380# 0.00133f
C1975 XA8.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C1976 D<6> XA1.XA3.MN0.G 0.0263f
C1977 XA0.XA6.MP0.G a_n232_47620# 4.4e-19
C1978 AVDD a_11000_42692# 0.358f
C1979 VREF a_22448_49028# 0.00255f
C1980 XA6.XA4.MN0.D a_14888_49028# 0.156f
C1981 AVDD a_9848_54308# 0.00166f
C1982 XA20.XA11.MN0.D XA20.XA11.MP0.D 0.0614f
C1983 a_8480_41636# a_8480_41284# 0.0109f
C1984 a_19928_41636# XA8.XA1.XA1.MN0.S 0.0674f
C1985 XA8.XA1.XA5.MN2.G XA7.XA1.XA2.MP0.D 0.146f
C1986 a_12368_47620# a_13520_47620# 0.00133f
C1987 XA4.XA4.MN0.G a_8480_46916# 2.84e-19
C1988 XA3.XA4.MN0.G a_9848_46916# 2.84e-19
C1989 AVDD a_7328_39876# 0.438f
C1990 XA3.XA4.MN0.D a_8480_45508# 9.24e-20
C1991 VREF a_12368_45508# 0.0556f
C1992 XA4.XA6.MP0.G SARP 0.0253f
C1993 XA0.XA7.MP0.G a_920_43396# 0.00442f
C1994 XA2.XA6.MP0.G a_5960_44452# 5.5e-19
C1995 XA2.XA11.MP0.D a_5960_52900# 0.00176f
C1996 AVDD a_2288_51844# 0.387f
C1997 XA5.XA11.MN1.G a_11000_52548# 9.29e-19
C1998 CK_SAMPLE SARN 0.00642f
C1999 a_7328_40228# a_7328_39876# 0.0109f
C2000 a_7328_45860# a_8480_45860# 0.00133f
C2001 XA1.XA4.MN0.G a_2288_43748# 6.3e-19
C2002 XA7.XA4.MN0.G XA7.XA1.XA5.MP1.D 0.00138f
C2003 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.D 0.0384f
C2004 XA6.XA1.XA5.MN2.G XA6.XA1.XA1.MP1.D 0.00107f
C2005 XA0.XA7.MP0.G a_n232_40932# 6.44e-19
C2006 XA4.XA6.MP0.G a_9848_42340# 7.76e-20
C2007 XA0.XA6.MP0.G a_n232_41988# 7.76e-20
C2008 XA4.XA9.MN1.G XA4.XA8.MP0.D 0.0132f
C2009 XA7.XA10.MP0.G XA8.XA1.XA5.MN2.G 2.18e-19
C2010 XA1.XA9.MN1.G a_2288_51492# 6.57e-19
C2011 a_18560_52196# XA7.XA7.MP0.D 0.0662f
C2012 AVDD a_23600_49732# 0.00154f
C2013 CK_SAMPLE a_9848_50084# 0.167f
C2014 XA8.XA9.MN1.G a_19928_51844# 0.0164f
C2015 a_13808_334# a_13808_n18# 0.0109f
C2016 XA1.XA4.MN0.D a_3440_40228# 4.11e-20
C2017 XA0.XA6.MP2.G XDAC1.XC0.XRES16.B 0.0333f
C2018 a_3440_44452# EN 0.00154f
C2019 a_920_44100# a_2288_44100# 8.89e-19
C2020 SARN li_14804_15696# 0.00103f
C2021 XA20.XA2a.MN0.D XA4.XA1.XA4.MP1.D 0.0128f
C2022 a_3440_45156# XA1.XA1.XA2.MP0.D 1.56e-20
C2023 D<5> a_7328_50788# 0.161f
C2024 a_11000_52196# VREF 0.00396f
C2025 XA2.XA1.XA5.MN2.G XA1.XA6.MP0.G 0.174f
C2026 AVDD a_920_46212# 0.356f
C2027 li_14804_19176# li_14804_18564# 0.00271f
C2028 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES8.B 0.0228f
C2029 XDAC2.XC128b<2>.XRES16.B XDAC2.XC128a<1>.XRES16.B 0.0114f
C2030 XA0.XA6.MP0.G XDAC2.XC64a<0>.XRES16.B 2.43e-19
C2031 a_920_43044# a_2288_43044# 8.89e-19
C2032 XA6.XA1.XA2.MP0.D XA6.XA1.XA4.MN1.D 0.056f
C2033 XA20.XA2a.MN0.D a_9848_40228# 2.1e-19
C2034 XA1.XA4.MN0.D XDAC1.XC128b<2>.XRES16.B 4.21e-20
C2035 XA0.XA4.MN0.D li_9184_20208# 0.00504f
C2036 AVDD XA7.XA1.XA5.MN0.D 0.00889f
C2037 XA8.XA7.MP0.G a_21080_47620# 0.00363f
C2038 a_14888_50084# XA6.XA4.MN0.D 3.12e-20
C2039 XA20.XA3.MN0.D a_23600_49732# 0.0585f
C2040 a_22448_50084# VREF 0.00119f
C2041 SARP a_9560_686# 2.97e-20
C2042 a_920_42340# XA0.XA1.XA1.MN0.S 1.34e-19
C2043 a_12368_41988# a_13520_41988# 0.00133f
C2044 XA2.XA6.MP0.G a_5960_45508# 5.5e-19
C2045 XA0.XA4.MN0.G a_920_47972# 0.155f
C2046 XA6.XA6.MP0.G a_16040_45860# 5.5e-19
C2047 XA20.XA9.MP0.D a_23600_42692# 0.14f
C2048 XA0.XA4.MN0.D a_920_46564# 2.2e-19
C2049 VREF a_n232_46564# 7.39e-19
C2050 AVDD XA6.XA1.XA1.MP1.D 0.0604f
C2051 XA6.XA1.XA5.MN2.G a_13520_44100# 2.31e-19
C2052 XA1.XA12.MP0.G a_3440_53252# 0.0661f
C2053 XA2.XA11.MN1.G a_4808_53252# 0.0689f
C2054 DONE a_23600_52900# 2.31e-19
C2055 a_9848_53604# a_11000_53604# 0.00133f
C2056 XA6.XA11.MN1.G XA5.XA11.MP0.D 0.0114f
C2057 AVDD XA20.XA4.MN0.D 0.456f
C2058 XA20.XA10.MN1.D a_23600_53604# 0.0269f
C2059 a_n232_40580# a_920_40580# 0.00133f
C2060 XA8.XA7.MP0.G a_21080_41988# 0.0719f
C2061 XA0.XA4.MN0.D XA0.XA1.XA5.MP0.D 9.69e-19
C2062 XA2.XA1.XA5.MN2.G a_4808_41636# 0.00417f
C2063 D<1> XA7.XA1.XA4.MP0.D 6.09e-19
C2064 D<5> a_8480_42340# 6.49e-19
C2065 XA5.XA6.MP0.G a_13520_43044# 7.76e-20
C2066 XA20.XA3.MN6.D a_22448_43396# 1.25e-19
C2067 XA0.XA11.MN1.G XB2.M1.G 0.22f
C2068 XA1.XA6.MP0.G XA1.XA1.XA4.MN1.D 7.41e-19
C2069 XA4.XA4.MN0.G a_9848_44804# 0.00858f
C2070 XA4.XA3.MN0.G a_9848_46212# 0.157f
C2071 XA0.XA10.MP0.G XA0.XA7.MP0.D 0.0601f
C2072 a_18560_52548# XA7.XA9.MN1.G 0.0711f
C2073 CK_SAMPLE a_8480_50788# 0.157f
C2074 a_5960_52548# a_5960_52196# 0.0109f
C2075 AVDD a_23600_50436# 0.00166f
C2076 XA2.XA9.MN1.G XA2.XA9.MN0.D 0.034f
C2077 a_8408_1742# a_9560_1742# 0.00133f
C2078 XA20.XA3a.MN0.D a_12368_42692# 0.00443f
C2079 XA5.XA6.MP0.G a_12368_40580# 5.5e-19
C2080 XA1.XA6.MP0.G a_2288_40228# 2.44e-19
C2081 XA0.XA4.MN0.G a_n232_42340# 7.97e-19
C2082 XA1.XA1.XA5.MN2.D a_2288_44100# 0.124f
C2083 a_3440_45508# EN 3.34e-19
C2084 a_5960_51140# a_7328_51140# 8.89e-19
C2085 XA8.XA1.XA5.MN2.G a_16040_51140# 7.1e-20
C2086 XA7.XA1.XA5.MN2.G a_17408_51140# 7.1e-20
C2087 AVDD a_n232_47268# 0.00125f
C2088 XA0.XA7.MP0.G XA0.XA6.MP2.G 0.624f
C2089 XA20.XA9.MP0.D XA8.XA4.MN0.D 0.0049f
C2090 XA3.XA7.MP0.D a_8480_50436# 1.37e-19
C2091 XB2.XA4.MP0.D XDAC2.XC1.XRES2.B 0.00369f
C2092 XA2.XA4.MN0.D XDAC1.XC0.XRES16.B 2.19e-20
C2093 EN a_22448_43044# 5.7e-20
C2094 XA20.XA2a.MN0.D a_18560_41284# 0.088f
C2095 XA4.XA1.XA2.MP0.D XA4.XA1.XA5.MP0.D 4.34e-19
C2096 D<1> XDAC1.XC32a<0>.XRES16.B 0.00136f
C2097 XA2.XA3.MN0.G a_4808_40932# 0.00369f
C2098 a_21080_50788# VREF 0.00361f
C2099 D<5> a_7328_49028# 0.00884f
C2100 AVDD a_13520_44100# 0.00125f
C2101 a_23600_50436# XA20.XA3.MN0.D 1.28e-19
C2102 D<1> a_17408_49380# 0.00891f
C2103 XA2.XA1.XA4.MN0.D a_5960_42340# 2.16e-19
C2104 XA2.XA1.XA4.MP0.D a_4808_42340# 2.16e-19
C2105 SARP a_22448_39876# 5.08e-19
C2106 D<8> li_14804_26136# 3.5e-20
C2107 EN a_21080_40580# 0.0714f
C2108 XA3.XA1.XA5.MN2.G a_5960_45156# 0.00486f
C2109 XA8.XA7.MP0.G XA8.XA1.XA5.MN2.D 0.108f
C2110 XA6.XA4.MN0.D a_16040_47972# 0.0546f
C2111 XA0.XA4.MN0.D XA20.XA3a.MN0.D 0.0705f
C2112 a_11000_48676# a_12368_48676# 8.89e-19
C2113 XA6.XA6.MP0.G a_14888_46916# 5e-19
C2114 XA3.XA6.MP0.G XA1.XA3.MN0.G 0.0276f
C2115 AVDD a_n232_41636# 0.00125f
C2116 XA0.XA6.MP0.G a_920_46564# 5.5e-19
C2117 D<3> a_14888_45860# 1.06e-19
C2118 AVDD a_22448_53604# 0.37f
C2119 a_2288_53956# XA2.XA11.MN1.G 0.0295f
C2120 a_16040_54308# XA7.XA11.MN1.G 0.00177f
C2121 XA6.XA1.XA1.MP2.D a_16040_40932# 0.00176f
C2122 a_16040_41284# XA6.XA1.XA1.MP1.D 0.00176f
C2123 a_4808_41284# a_4808_40932# 0.0109f
C2124 XA3.XA4.MN0.G a_9848_45860# 2.2e-19
C2125 XA4.XA4.MN0.G a_8480_45860# 2.2e-19
C2126 AVDD a_8408_1390# 0.435f
C2127 a_5960_46916# a_7328_46916# 8.89e-19
C2128 XA5.XA1.XA5.MN2.G a_11000_42692# 0.00442f
C2129 VREF a_11000_44452# 0.0182f
C2130 XA3.XA4.MN0.D a_7328_44452# 9.15e-20
C2131 XA0.XA6.MP0.G XA0.XA1.XA5.MP0.D 0.00121f
C2132 a_4808_52900# a_4808_52548# 0.0109f
C2133 a_14888_52900# XA6.XA10.MP0.G 0.0681f
C2134 XA6.XA10.MP0.D a_14888_52548# 0.00316f
C2135 AVDD a_18560_51140# 0.00166f
C2136 CK_SAMPLE a_14888_51492# 6.34e-19
C2137 XA5.XA11.MN1.G a_13520_51844# 3.12e-19
C2138 a_8408_3502# XB1.XA1.MP0.D 1.47e-19
C2139 D<4> a_11000_40580# 4.07e-20
C2140 XA4.XA1.XA5.MN2.G a_8480_39876# 2.97e-20
C2141 XA0.XA6.MP2.G a_920_40228# 7.76e-20
C2142 XA7.XA3.MN0.G a_18560_44100# 0.00441f
C2143 XA2.XA3.MN0.G EN 0.0863f
C2144 XA20.XA3a.MN0.D XA8.XA1.XA2.MP0.D 0.193f
C2145 XA1.XA1.XA5.MN2.D XA2.XA1.XA5.MN2.D 0.00869f
C2146 a_8480_45508# a_8480_45156# 0.0109f
C2147 XA6.XA6.MP0.G XA6.XA1.XA1.MN0.S 0.0173f
C2148 XA2.XA4.MN0.G a_4808_43044# 0.0409f
C2149 XA7.XA12.MP0.G VREF 0.0123f
C2150 XA20.XA10.MN1.D a_23600_49732# 0.00444f
C2151 XA2.XA8.MP0.D a_4808_51492# 0.00224f
C2152 a_16040_51844# a_16040_51492# 0.0109f
C2153 XA5.XA9.MN1.G D<3> 0.0378f
C2154 AVDD a_23600_48676# 0.00154f
C2155 CK_SAMPLE a_8480_49028# 7.31e-19
C2156 XA2.XA7.MP0.D a_4808_51140# 0.00388f
C2157 XA20.XA4.MN0.D a_23600_50788# 0.0584f
C2158 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES2.B 0.0136f
C2159 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES8.B 0.471f
C2160 XA20.XA3a.MN0.D XA7.XA1.XA1.MP1.D 0.0093f
C2161 XA0.XA6.MP2.G li_9184_20820# 3.5e-20
C2162 XA3.XA1.XA5.MP1.D a_8480_43748# 2.16e-19
C2163 XA3.XA1.XA5.MN1.D a_7328_43748# 2.16e-19
C2164 XA20.XA2a.MN0.D a_2288_41988# 0.00302f
C2165 XA3.XA3.MN0.G a_9848_41636# 7.98e-19
C2166 EN a_17408_43748# 0.166f
C2167 a_21080_44100# a_21080_43748# 0.0109f
C2168 AVDD a_2288_45156# 0.356f
C2169 XA3.XA1.XA5.MN2.G VREF 0.704f
C2170 XA2.XA1.XA5.MN2.G XA1.XA4.MN0.D 0.198f
C2171 a_23600_50788# a_23600_50436# 0.0109f
C2172 D<5> a_7328_50084# 0.0155f
C2173 XDAC1.XC32a<0>.XRES4.B XDAC1.XC64a<0>.XRES4.B 0.00284f
C2174 li_9184_13860# li_9184_13248# 0.00271f
C2175 XA0.XA4.MN0.D XDAC1.XC64a<0>.XRES16.B 2.43e-19
C2176 XA1.XA4.MN0.D li_9184_10380# 0.00504f
C2177 XA8.XA1.XA4.MN1.D XA8.XA1.XA4.MP1.D 0.00918f
C2178 D<3> a_13520_46916# 0.00249f
C2179 XA4.XA6.MP0.G a_9848_47972# 6.28e-19
C2180 a_4808_49380# a_4808_49028# 0.0109f
C2181 XA8.XA7.MP0.G a_22448_46564# 8.22e-19
C2182 XA7.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.51f
C2183 D<7> XA3.XA3.MN0.G 0.16f
C2184 D<6> D<8> 0.0323f
C2185 XA0.XA6.MP0.G XA20.XA3a.MN0.D 0.0687f
C2186 AVDD a_9848_42692# 0.00125f
C2187 XA20.XA3.MN0.D a_23600_48676# 0.0297f
C2188 VREF a_21080_49028# 0.0646f
C2189 AVDD a_8480_54308# 0.00166f
C2190 XA20.XA11.MN0.D DONE 0.12f
C2191 SARP XDAC1.X16ab.XRES4.B 13.9f
C2192 D<1> XA7.XA1.XA5.MN1.D 0.00185f
C2193 XA7.XA1.XA5.MN2.G XA7.XA1.XA2.MP0.D 0.126f
C2194 XA3.XA4.MN0.G a_8480_46916# 0.0885f
C2195 AVDD a_5960_39876# 0.44f
C2196 XA3.XA4.MN0.D a_7328_45508# 9.15e-20
C2197 VREF a_11000_45508# 0.0556f
C2198 XA0.XA7.MP0.G a_n232_43396# 1.95e-19
C2199 XA2.XA6.MP0.G a_4808_44452# 7.76e-20
C2200 a_n232_47620# a_n232_47268# 0.0109f
C2201 XA6.XA6.MP0.G a_16040_44804# 5.5e-19
C2202 a_16040_53252# a_17408_53252# 8.89e-19
C2203 a_5960_53252# XA2.XA10.MP0.D 0.0661f
C2204 XA8.XA11.MP0.D XA8.XA10.MP0.D 0.00986f
C2205 XA20.XA10.MN1.D XA20.XA4.MN0.D 0.11f
C2206 AVDD a_920_51844# 0.387f
C2207 CK_SAMPLE XA8.XA9.MN0.D 1.12e-19
C2208 a_9848_53956# XA4.XA9.MN1.G 7.37e-20
C2209 a_18560_40228# a_19928_40228# 8.89e-19
C2210 a_19928_46212# a_19928_45860# 0.0109f
C2211 XA4.XA3.MN0.G a_11000_45156# 0.0546f
C2212 XA6.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.D 0.0288f
C2213 XA1.XA4.MN0.D XA1.XA1.XA4.MN1.D 9.89e-19
C2214 a_2288_52548# XA2.XA1.XA5.MN2.G 1.75e-19
C2215 a_17408_52196# XA7.XA7.MP0.D 0.0674f
C2216 XA0.XA7.MP0.D XA1.XA7.MP0.D 0.00435f
C2217 AVDD a_22448_49732# 0.417f
C2218 CK_SAMPLE a_8480_50084# 0.167f
C2219 XA20.XA10.MN1.D a_23600_50436# 0.0744f
C2220 a_7328_52196# a_7328_51844# 0.0109f
C2221 XA8.XA9.MN1.G a_18560_51844# 2.2e-19
C2222 a_8408_n18# a_9560_n18# 0.00133f
C2223 a_2288_44452# EN 0.00173f
C2224 a_13520_44452# a_13520_44100# 0.0109f
C2225 XA1.XA4.MN0.D a_2288_40228# 4.07e-20
C2226 XA20.XA2a.MN0.D XA4.XA1.XA4.MN1.D 0.0128f
C2227 XA0.XA7.MP0.G XA1.XA6.MP0.G 0.0666f
C2228 AVDD a_n232_46212# 0.00125f
C2229 a_21080_51140# a_21080_50788# 0.0109f
C2230 a_13520_43396# a_13520_43044# 0.0109f
C2231 XA2.XA1.XA2.MP0.D a_5960_42692# 7.68e-20
C2232 XA20.XA2a.MN0.D a_8480_40228# 2.1e-19
C2233 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES2.B 0.00405f
C2234 AVDD XA7.XA1.XA5.MP0.D 0.159f
C2235 D<5> a_8480_47972# 5.43e-19
C2236 a_21080_50084# VREF 0.00526f
C2237 a_23600_50084# a_23600_49732# 0.0109f
C2238 a_9848_49732# a_11000_49732# 0.00133f
C2239 a_n232_41988# a_n232_41636# 0.0109f
C2240 a_12368_48324# a_12368_47972# 0.0109f
C2241 XA6.XA6.MP0.G a_14888_45860# 1.38e-19
C2242 XA4.XA4.MN0.G XA5.XA4.MN0.G 0.00869f
C2243 XA0.XA4.MN0.G a_n232_47972# 0.153f
C2244 D<7> a_3440_44452# 5.26e-19
C2245 XA20.XA9.MP0.D a_22448_42692# 0.066f
C2246 XA0.XA4.MN0.D a_n232_46564# 0.001f
C2247 AVDD XA6.XA1.XA1.MN0.D 0.0357f
C2248 XA4.XA4.MN0.D XA4.XA3.MN0.G 0.00642f
C2249 VREF XA8.XA3.MN0.G 0.603f
C2250 XA5.XA1.XA5.MN2.G a_13520_44100# 0.0693f
C2251 XA6.XA1.XA5.MN2.G a_12368_44100# 0.00556f
C2252 XA2.XA6.MP0.G a_4808_45508# 7.76e-20
C2253 XA2.XA11.MN1.G a_3440_53252# 0.0238f
C2254 XA1.XA12.MP0.G a_2288_53252# 0.00276f
C2255 AVDD XA8.XA10.MP0.G 0.855f
C2256 XA20.XA10.MN1.D a_22448_53604# 0.0448f
C2257 XA20.XA11.MN0.D a_23600_52900# 1.46e-19
C2258 DONE a_22448_52900# 0.00597f
C2259 a_12368_40932# a_12368_40580# 0.0109f
C2260 XA8.XA7.MP0.G a_19928_41988# 0.0684f
C2261 XA0.XA4.MN0.D XA0.XA1.XA5.MN0.D 9.9e-19
C2262 XA2.XA1.XA5.MN2.G a_3440_41636# 0.131f
C2263 XA0.XA11.MN1.G XB1.XA4.MN0.D 7.05e-19
C2264 D<5> a_7328_42340# 7.77e-20
C2265 XA5.XA6.MP0.G a_12368_43044# 5.5e-19
C2266 XA20.XA3a.MN0.G a_22448_43396# 1.63e-19
C2267 a_13520_46564# a_14888_46564# 8.89e-19
C2268 a_920_46564# a_920_46212# 0.0109f
C2269 XA1.XA6.MP0.G XA1.XA1.XA4.MP1.D 0.00121f
C2270 XA3.XA4.MN0.G a_9848_44804# 2.2e-19
C2271 XA4.XA4.MN0.G a_8480_44804# 2.2e-19
C2272 XA6.XA10.MP0.G a_16040_52196# 0.0441f
C2273 a_17408_52548# XA7.XA9.MN1.G 0.0674f
C2274 CK_SAMPLE a_7328_50788# 0.00142f
C2275 AVDD a_22448_50436# 0.389f
C2276 XB2.XA4.MP0.D XB2.XA3.MN1.D 0.376p
C2277 SAR_IP a_11000_686# 0.0598f
C2278 a_13808_2094# a_13808_1742# 0.0109f
C2279 XA20.XA3a.MN0.D a_11000_42692# 0.00443f
C2280 a_21080_45156# a_21080_44804# 0.0109f
C2281 a_7328_44804# a_8480_44804# 0.00133f
C2282 XA6.XA4.MN0.G XA6.XA1.XA4.MN0.D 0.00331f
C2283 XA2.XA3.MN0.G a_4808_43396# 0.00341f
C2284 XA7.XA1.XA5.MN2.D a_18560_44452# 0.153f
C2285 a_2288_45508# EN 1.42e-19
C2286 XA3.XA4.MN0.D a_8480_41284# 9.24e-20
C2287 SARN li_14804_26136# 0.00103f
C2288 XA20.XA10.MN1.D a_23600_48676# 0.00405f
C2289 XA7.XA1.XA5.MN2.G a_16040_51140# 0.077f
C2290 AVDD a_23600_47620# 0.00154f
C2291 a_7328_52900# VREF 0.00396f
C2292 XB1.XA4.MP0.D XDAC1.XC1.XRES16.B 0.0646f
C2293 li_14804_24300# li_14804_23688# 0.00271f
C2294 XDAC2.X16ab.XRES2.B XDAC2.X16ab.XRES1A.B 0.0136f
C2295 XDAC1.X16ab.XRES16.B li_9184_23688# 0.00117f
C2296 XDAC2.X16ab.XRES4.B XDAC2.XC128b<2>.XRES4.B 0.00284f
C2297 EN a_21080_43044# 0.14f
C2298 XA1.XA4.MN0.D XDAC1.XC0.XRES16.B 4.21e-20
C2299 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES16.B 0.0301f
C2300 XA20.XA2a.MN0.D a_17408_41284# 0.0685f
C2301 XA4.XA1.XA2.MP0.D XA4.XA1.XA5.MN0.D 0.056f
C2302 a_11000_43748# a_11000_43396# 0.0109f
C2303 XA1.XA3.MN0.G a_4808_40932# 4.4e-20
C2304 XA2.XA3.MN0.G a_3440_40932# 4.21e-19
C2305 AVDD a_12368_44100# 0.359f
C2306 XA3.XA6.MN0.D a_8480_50084# 0.0488f
C2307 a_23600_50436# a_23600_50084# 0.0109f
C2308 XA2.XA1.XA5.MN2.G a_2288_48324# 0.00455f
C2309 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES4.B 0.428f
C2310 a_17408_42692# a_17408_42340# 0.0109f
C2311 XA2.XA1.XA4.MN0.D a_4808_42340# 0.0474f
C2312 XA7.XA1.XA2.MP0.D a_17408_41284# 1.07e-19
C2313 XA3.XA1.XA5.MN2.G a_4808_45156# 1.95e-19
C2314 XA8.XA1.XA5.MN2.G XA8.XA1.XA5.MN2.D 0.0398f
C2315 D<7> a_3440_45508# 0.0031f
C2316 XA6.XA4.MN0.D a_14888_47972# 0.0788f
C2317 VREF a_22448_47972# 0.00191f
C2318 a_23600_49028# a_23600_48676# 0.0109f
C2319 AVDD a_23600_41988# 0.00193f
C2320 XA20.XA3.MN0.D a_23600_47620# 0.0276f
C2321 XA0.XA6.MP0.G a_n232_46564# 7.76e-20
C2322 XA2.XA6.MP0.G XA3.XA3.MN0.G 3.56f
C2323 D<3> a_13520_45860# 0.0675f
C2324 XA3.XA6.MP0.G D<8> 0.0791f
C2325 a_13520_53956# a_14888_53956# 8.89e-19
C2326 a_3440_53956# XA0.XA12.MP0.D 0.00258f
C2327 AVDD a_21080_53604# 0.384f
C2328 a_14888_54308# XA7.XA11.MN1.G 2.54e-19
C2329 XA1.XA1.XA1.MN0.S a_3440_40580# 0.00155f
C2330 XA6.XA1.XA1.MN0.S a_16040_40932# 0.0271f
C2331 SARP li_9184_15696# 0.00103f
C2332 XA3.XA4.MN0.G a_8480_45860# 0.0146f
C2333 AVDD XB2.XA3.MN1.D 1.65f
C2334 a_8480_47268# XA3.XA3.MN0.G 2.69e-19
C2335 a_18560_47268# a_18560_46916# 0.0109f
C2336 XA0.XA6.MP2.G XA0.XA1.XA4.MP1.D 7.42e-19
C2337 XA4.XA1.XA5.MN2.G a_11000_42692# 1.97e-19
C2338 XA5.XA1.XA5.MN2.G a_9848_42692# 1.95e-19
C2339 D<4> a_11000_43044# 7.76e-20
C2340 XA4.XA6.MP0.G a_11000_43748# 5.5e-19
C2341 VREF a_9848_44452# 7.12e-19
C2342 XA0.XA6.MP0.G XA0.XA1.XA5.MN0.D 7.41e-19
C2343 a_22448_52900# a_23600_52900# 0.00133f
C2344 AVDD a_17408_51140# 0.383f
C2345 CK_SAMPLE a_13520_51492# 6.45e-19
C2346 XA5.XA11.MN1.G a_12368_51844# 4.48e-19
C2347 a_9560_3854# XB1.XA1.MP0.D 1.01e-19
C2348 a_9560_3150# a_9560_2798# 0.0109f
C2349 a_13808_3502# a_13808_3150# 0.0109f
C2350 a_14960_3502# XB2.XA2.MN0.G 0.0939f
C2351 D<4> a_9848_40580# 5.24e-19
C2352 XA3.XA1.XA5.MN2.G a_8480_39876# 0.00325f
C2353 XA4.XA1.XA5.MN2.G a_7328_39876# 8.8e-19
C2354 XA0.XA6.MP2.G a_n232_40228# 6.49e-19
C2355 XA7.XA3.MN0.G a_17408_44100# 0.00245f
C2356 XA1.XA3.MN0.G EN 0.0841f
C2357 D<8> XA0.XA1.XA5.MN1.D 8.47e-19
C2358 XA20.XA3.MN0.D a_23600_41988# 8.5e-20
C2359 XA2.XA6.MP0.G a_5960_41284# 4.24e-19
C2360 XA20.XA3a.MN0.D XA7.XA1.XA5.MN0.D 0.0111f
C2361 a_18560_45508# XA7.XA1.XA5.MN2.D 0.0658f
C2362 XA8.XA4.MN0.G a_21080_43396# 8.07e-19
C2363 XA20.XA10.MN1.D a_22448_49732# 1.87e-19
C2364 XA8.XA11.MN1.G VREF 0.017f
C2365 SARN D<6> 0.027f
C2366 a_2288_52196# D<7> 7.56e-20
C2367 AVDD a_22448_48676# 0.438f
C2368 CK_SAMPLE a_7328_49028# 3.27e-19
C2369 XA20.XA4.MN0.D a_22448_50788# 0.00246f
C2370 XA7.XA7.MP0.D XA8.XA1.XA5.MN2.G 0.14f
C2371 XA20.XA3a.MN0.D XA6.XA1.XA1.MP1.D 0.0093f
C2372 XA3.XA1.XA5.MP1.D a_7328_43748# 0.049f
C2373 XA20.XA2a.MN0.D a_920_41988# 0.00302f
C2374 XA3.XA3.MN0.G a_8480_41636# 0.00333f
C2375 EN a_16040_43748# 0.166f
C2376 a_9848_50436# a_11000_50436# 0.00133f
C2377 AVDD a_920_45156# 0.356f
C2378 XA0.XA7.MP0.G XA1.XA4.MN0.D 0.069f
C2379 XA2.XA1.XA5.MN2.G VREF 0.704f
C2380 D<1> XA7.XA6.MN0.D 0.00148f
C2381 XA3.XA1.XA4.MN1.D a_8480_42692# 0.0474f
C2382 a_21080_43044# a_21080_42692# 0.0109f
C2383 XA20.XA3.MN1.D a_23600_48324# 0.00245f
C2384 D<3> a_12368_46916# 0.0185f
C2385 a_16040_49380# a_17408_49380# 8.89e-19
C2386 XA8.XA7.MP0.G a_21080_46564# 0.00363f
C2387 XA6.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C2388 D<7> XA2.XA3.MN0.G 0.112f
C2389 AVDD a_8480_42692# 0.00125f
C2390 XA7.XA6.MP0.G XA7.XA4.MN0.G 0.0415f
C2391 XA5.XA4.MN0.D a_13520_49028# 0.156f
C2392 VREF a_19928_49028# 7.81e-19
C2393 XA20.XA9.MP0.D EN 0.00951f
C2394 AVDD a_7328_54308# 0.448f
C2395 a_23600_54660# DONE 0.0658f
C2396 a_22448_54660# XA20.XA11.MP0.D 0.00176f
C2397 a_7328_41636# a_7328_41284# 0.0109f
C2398 XA2.XA1.XA1.MN0.S XA3.XA1.XA1.MN0.S 0.00217f
C2399 D<1> XA7.XA1.XA5.MP1.D 7.43e-19
C2400 XA7.XA1.XA5.MN2.G XA6.XA1.XA5.MP0.D 0.00353f
C2401 a_11000_47620# a_12368_47620# 8.89e-19
C2402 XA3.XA4.MN0.G a_7328_46916# 0.0662f
C2403 AVDD a_4808_39876# 0.00131f
C2404 SARN a_23600_42692# 0.00204f
C2405 XA6.XA6.MP0.G a_14888_44804# 7.76e-20
C2406 a_4808_53252# XA2.XA10.MP0.D 0.0692f
C2407 AVDD a_n232_51844# 0.00166f
C2408 DONE a_23600_52196# 1.97e-19
C2409 CK_SAMPLE XA8.XA9.MN1.G 0.193f
C2410 a_5960_40228# a_5960_39876# 0.0109f
C2411 D<3> XA5.XA1.XA1.MN0.S 0.0157f
C2412 a_5960_45860# a_7328_45860# 8.89e-19
C2413 XA0.XA4.MN0.G a_920_43748# 6.3e-19
C2414 XA4.XA3.MN0.G a_9848_45156# 0.0805f
C2415 XA6.XA4.MN0.G XA6.XA1.XA5.MP1.D 0.00138f
C2416 XA20.XA3a.MN0.D a_13520_44100# 5.04e-20
C2417 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.D 0.0825f
C2418 XA1.XA4.MN0.D XA1.XA1.XA4.MP1.D 9.71e-19
C2419 XA6.XA10.MP0.G XA7.XA1.XA5.MN2.G 2.18e-19
C2420 XA7.XA9.MN0.D a_18560_51844# 0.00176f
C2421 XA7.XA9.MN1.G a_19928_51844# 2.2e-19
C2422 AVDD a_21080_49732# 0.36f
C2423 CK_SAMPLE a_7328_50084# 0.00848f
C2424 XA20.XA10.MN1.D a_22448_50436# 0.0658f
C2425 a_12368_334# a_12368_n18# 0.0109f
C2426 XA0.XA6.MP2.G li_9184_31260# 0.00508f
C2427 a_920_44452# EN 0.00173f
C2428 a_n232_44100# a_920_44100# 0.00133f
C2429 XA20.XA3a.MN0.D a_n232_41636# 0.00542f
C2430 SARN XDAC2.XC32a<0>.XRES1B.B 3.59f
C2431 XA20.XA2a.MN0.D XA3.XA1.XA4.MN1.D 0.0128f
C2432 XA3.XA4.MN0.G XA3.XA1.XA1.MN0.S 5.22e-20
C2433 XA4.XA9.MN1.G a_11000_49380# 2.54e-19
C2434 AVDD XA20.XA2a.MN0.D 9.22f
C2435 XA20.XA10.MN1.D a_23600_47620# 0.00423f
C2436 XA2.XA6.MP2.D a_5960_50788# 0.049f
C2437 li_9184_19176# li_9184_18564# 0.00271f
C2438 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES8.B 0.0228f
C2439 XDAC1.XC128b<2>.XRES16.B XDAC1.XC128a<1>.XRES16.B 0.0114f
C2440 XA0.XA6.MP0.G li_14804_10380# 1.85e-20
C2441 a_n232_43044# a_920_43044# 0.00133f
C2442 XA2.XA1.XA2.MP0.D a_4808_42692# 0.0962f
C2443 XA0.XA4.MN0.D XDAC1.XC128b<2>.XRES16.B 0.0301f
C2444 EN a_12368_42340# 0.159f
C2445 XA2.XA1.XA5.MN2.G a_2288_47268# 0.00363f
C2446 AVDD XA7.XA1.XA2.MP0.D 0.263f
C2447 D<5> a_7328_47972# 0.0147f
C2448 D<2> XA6.XA4.MN0.G 0.26f
C2449 a_13520_50084# XA5.XA4.MN0.D 3.12e-20
C2450 a_11000_41988# a_12368_41988# 8.89e-19
C2451 D<3> a_13520_44804# 5.26e-19
C2452 D<7> a_2288_44452# 1.48e-19
C2453 D<6> SARP 0.0759f
C2454 XA20.XA10.MN1.D a_23600_41988# 0.00492f
C2455 XA20.XA3.MN0.D XA20.XA2a.MN0.D 0.218f
C2456 AVDD XA5.XA1.XA1.MN0.D 0.0357f
C2457 VREF XA7.XA3.MN0.G 0.608f
C2458 XA5.XA1.XA5.MN2.G a_12368_44100# 7.1e-20
C2459 XA6.XA1.XA5.MN2.G a_11000_44100# 7.1e-20
C2460 XA2.XA11.MN1.G a_2288_53252# 3.16e-19
C2461 a_8480_53604# a_9848_53604# 8.89e-19
C2462 AVDD XA7.XA10.MP0.G 0.853f
C2463 XA0.XA12.MP0.D a_4808_53252# 2.81e-19
C2464 XA5.XA11.MN1.G XA5.XA11.MP0.D 0.0383f
C2465 XA4.XA12.MP0.G XA4.XA11.MP0.D 0.0612f
C2466 DONE a_21080_52900# 0.00176f
C2467 XA8.XA1.XA5.MN2.G a_19928_41988# 0.00407f
C2468 XA0.XA4.MN0.D XA0.XA1.XA2.MP0.D 0.0111f
C2469 XA2.XA1.XA5.MN2.G a_2288_41636# 0.0736f
C2470 XA0.XA7.MP0.G a_3440_41636# 0.0039f
C2471 XA0.XA11.MN1.G XB1.XA4.MP0.D 7.2e-20
C2472 XA3.XA4.MN0.G a_8480_44804# 0.00858f
C2473 XA3.XA3.MN0.G a_8480_46212# 0.157f
C2474 CK_SAMPLE a_5960_50788# 0.00142f
C2475 a_4808_52548# a_4808_52196# 0.0109f
C2476 XA6.XA10.MP0.G a_14888_52196# 0.0131f
C2477 AVDD a_21080_50436# 0.417f
C2478 XB2.XA4.MP0.D XB2.XA3.MN0.S 1.67e-19
C2479 a_8408_2094# XB1.XA3.MN1.D 0.00291f
C2480 SAR_IP a_9560_686# 5.55e-19
C2481 XB1.XA0.MP0.D a_9560_1742# 0.0797f
C2482 a_9560_2094# XB1.XA3.MN0.S 3.29e-19
C2483 XA20.XA3a.MN0.D a_9848_42692# 0.0099f
C2484 XA20.XA2a.MN0.D XA1.XA1.XA2.MP0.D 0.227f
C2485 XA8.XA3.MN0.G XA8.XA1.XA2.MP0.D 0.00212f
C2486 XA1.XA3.MN0.G a_4808_43396# 4.4e-20
C2487 XA2.XA3.MN0.G a_3440_43396# 4.21e-19
C2488 XA0.XA1.XA5.MN2.D a_920_44100# 0.126f
C2489 XA7.XA1.XA5.MN2.D a_17408_44452# 0.158f
C2490 a_920_45508# EN 1.42e-19
C2491 XA3.XA4.MN0.D a_7328_41284# 9.15e-20
C2492 XA7.XA1.XA5.MN2.G a_14888_51140# 0.0661f
C2493 a_4808_51140# a_5960_51140# 0.00133f
C2494 XA20.XA10.MN1.D a_22448_48676# 1.78e-19
C2495 AVDD a_22448_47620# 0.369f
C2496 a_23600_51492# a_23600_51140# 0.0109f
C2497 SARN XA3.XA6.MP0.G 0.0424f
C2498 XA20.XA4.MN0.D a_22448_50084# 2.11e-19
C2499 a_5960_52900# VREF 0.00396f
C2500 XA5.XA9.MN1.G XA5.XA6.MN0.D 0.0615f
C2501 EN a_19928_43044# 1.25e-19
C2502 XA20.XA2a.MN0.D a_16040_41284# 0.0669f
C2503 SARP a_23600_42692# 0.02f
C2504 XA1.XA3.MN0.G a_3440_40932# 0.00366f
C2505 AVDD a_11000_44100# 0.359f
C2506 XA0.XA7.MP0.G a_2288_48324# 7.1e-20
C2507 XA2.XA1.XA5.MN2.G a_920_48324# 7.1e-20
C2508 D<8> XDAC2.X16ab.XRES1B.B 4.06e-21
C2509 XA8.XA1.XA5.MN2.G XA7.XA1.XA5.MN2.D 0.108f
C2510 D<7> a_2288_45508# 0.00436f
C2511 VREF a_21080_47972# 0.0171f
C2512 AVDD a_22448_41988# 0.57f
C2513 XA2.XA1.XA5.MN2.G a_4808_45156# 1e-19
C2514 XA2.XA6.MP0.G XA2.XA3.MN0.G 3.15f
C2515 D<3> a_12368_45860# 0.0774f
C2516 a_9848_48676# a_11000_48676# 0.00133f
C2517 a_2288_53956# XA0.XA12.MP0.D 0.00198f
C2518 a_920_53956# XA0.XA12.MP0.G 0.0658f
C2519 AVDD a_19928_53604# 0.00166f
C2520 XA1.XA1.XA1.MN0.S a_2288_40580# 0.0318f
C2521 a_14888_41284# XA6.XA1.XA1.MN0.D 0.00224f
C2522 a_3440_41284# a_3440_40932# 0.0109f
C2523 XA3.XA4.MN0.G a_7328_45860# 2.12e-19
C2524 AVDD XB2.XA3.MN0.S 0.183f
C2525 a_4808_46916# a_5960_46916# 0.00133f
C2526 XA0.XA6.MP2.G XA0.XA1.XA4.MN1.D 0.00188f
C2527 XA4.XA1.XA5.MN2.G a_9848_42692# 0.0739f
C2528 D<4> a_9848_43044# 6.49e-19
C2529 XA4.XA6.MP0.G a_9848_43748# 7.76e-20
C2530 XA2.XA4.MN0.D a_5960_44452# 9.14e-20
C2531 VREF a_8480_44452# 7.12e-19
C2532 XA0.XA6.MP0.G XA0.XA1.XA2.MP0.D 0.0106f
C2533 a_9848_53252# XA4.XA9.MN1.G 5.25e-19
C2534 a_3440_52900# a_3440_52548# 0.0109f
C2535 a_13520_52900# XA5.XA10.MP0.G 0.0665f
C2536 XA5.XA10.MP0.D a_13520_52548# 0.00316f
C2537 AVDD a_16040_51140# 0.383f
C2538 CK_SAMPLE a_12368_51492# 5.02e-19
C2539 XA5.XA11.MN1.G a_11000_51844# 2.62e-19
C2540 a_8408_3854# XB1.XA1.MP0.D 7.02e-20
C2541 a_13808_3502# XB2.XA2.MN0.G 0.0674f
C2542 XA3.XA1.XA5.MN2.G a_7328_39876# 0.00278f
C2543 D<8> EN 0.298f
C2544 SARN a_13808_1038# 2.97e-20
C2545 XA2.XA6.MP0.G a_4808_41284# 3.97e-20
C2546 XA20.XA3a.MN0.D XA7.XA1.XA5.MP0.D 7.25e-19
C2547 XA0.XA1.XA5.MN2.D XA1.XA1.XA5.MN2.D 0.00869f
C2548 a_17408_45508# XA7.XA1.XA5.MN2.D 0.0675f
C2549 a_7328_45508# a_7328_45156# 0.0109f
C2550 XA6.XA6.MP0.G XA5.XA1.XA1.MN0.S 4.2e-19
C2551 XA1.XA4.MN0.G a_3440_43044# 0.0409f
C2552 XA8.XA4.MN0.G a_19928_43396# 0.0104f
C2553 XA1.XA8.MP0.D a_3440_51492# 0.00224f
C2554 a_14888_51844# a_14888_51492# 0.0109f
C2555 XA6.XA12.MP0.G VREF 0.0119f
C2556 AVDD a_21080_48676# 0.356f
C2557 CK_SAMPLE a_5960_49028# 3.27e-19
C2558 XA1.XA7.MP0.D a_3440_51140# 0.00388f
C2559 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES8.B 0.0228f
C2560 XDAC2.XC0.XRES16.B XDAC2.XC64b<1>.XRES16.B 0.0114f
C2561 li_14804_29616# li_14804_29004# 0.00271f
C2562 XA20.XA3a.MN0.D XA6.XA1.XA1.MN0.D 0.0616f
C2563 XA0.XA6.MP2.G XDAC1.XC128b<2>.XRES2.B 4.06e-21
C2564 XA7.XA1.XA5.MP1.D XA7.XA1.XA5.MN1.D 0.00918f
C2565 XA20.XA2a.MN0.D a_n232_41988# 0.0844f
C2566 SARN li_14804_5676# 0.00228f
C2567 EN a_14888_43748# 0.00532f
C2568 a_19928_44100# a_19928_43748# 0.0109f
C2569 XA0.XA6.MP0.G XDAC2.XC0.XRES16.B 8.44e-20
C2570 XA20.XA10.MN1.D XA20.XA2a.MN0.D 0.0217f
C2571 AVDD a_n232_45156# 0.00125f
C2572 a_8480_50788# XA3.XA6.MP0.G 1.75e-20
C2573 XA8.XA1.XA5.MN2.G a_17408_49732# 0.00457f
C2574 D<1> XA7.XA6.MP0.D 0.0323f
C2575 XA2.XA1.XA5.MN2.G XA0.XA4.MN0.D 6.95e-19
C2576 XA0.XA7.MP0.G VREF 0.704f
C2577 a_22448_50788# a_22448_50436# 0.0109f
C2578 XDAC2.XC32a<0>.XRES2.B XDAC2.XC32a<0>.XRES16.B 0.457f
C2579 EN a_2288_41284# 0.00564f
C2580 XA0.XA4.MN0.D li_9184_10380# 1.85e-20
C2581 XA1.XA4.MN0.D XDAC1.XC64a<0>.XRES2.B 0.00405f
C2582 XA8.XA1.XA2.MP0.D a_21080_42340# 2.54e-19
C2583 XA3.XA1.XA4.MN1.D a_7328_42692# 2.16e-19
C2584 XA3.XA1.XA4.MP1.D a_8480_42692# 2.16e-19
C2585 XA0.XA1.XA2.MP0.D a_920_41636# 0.00224f
C2586 XA4.XA1.XA2.MP0.D a_11000_41988# 0.0219f
C2587 XA20.XA3.MN6.D a_23600_48324# 5.76e-19
C2588 XA20.XA3.MN1.D a_22448_48324# 0.00245f
C2589 XA5.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.51f
C2590 XA2.XA1.XA5.MN2.G a_2288_46212# 0.00363f
C2591 D<7> XA1.XA3.MN0.G 1.21f
C2592 AVDD a_7328_42692# 0.358f
C2593 XA5.XA4.MN0.D a_12368_49028# 0.154f
C2594 a_3440_49380# a_3440_49028# 0.0109f
C2595 VREF a_18560_49028# 7.81e-19
C2596 XA20.XA9.MP0.D a_23600_44100# 0.00334f
C2597 AVDD a_5960_54308# 0.447f
C2598 a_23600_54660# XA20.XA11.MN0.D 0.00437f
C2599 a_22448_54660# DONE 0.0714f
C2600 XA20.XA12.MP0.G XA20.XA11.MP0.D 0.00409f
C2601 a_17408_41636# XA7.XA1.XA1.MP2.D 0.00176f
C2602 a_18560_41636# XA7.XA1.XA1.MN0.S 0.0658f
C2603 XA2.XA1.XA1.MN0.S XA2.XA1.XA1.MP2.D 0.0708f
C2604 SARP li_9184_26136# 0.00103f
C2605 XA7.XA1.XA5.MN2.G XA6.XA1.XA5.MN0.D 7.2e-19
C2606 AVDD a_3440_39876# 0.00131f
C2607 XA2.XA4.MN0.D a_5960_45508# 9.14e-20
C2608 D<5> a_8480_43748# 6.49e-19
C2609 XA20.XA3a.MN0.D a_23600_47620# 0.0526f
C2610 XA3.XA6.MP0.G SARP 0.0253f
C2611 XA4.XA11.MN1.G a_9848_52548# 2.85e-19
C2612 AVDD XA8.XA7.MP0.D 1.2f
C2613 DONE a_22448_52196# 0.00486f
C2614 XA7.XA11.MP0.D XA7.XA10.MP0.D 0.00986f
C2615 a_14888_53252# a_16040_53252# 0.00133f
C2616 a_17408_40228# a_18560_40228# 0.00133f
C2617 a_18560_46212# a_18560_45860# 0.0109f
C2618 XA6.XA4.MN0.G XA6.XA1.XA5.MN1.D 0.0242f
C2619 XA0.XA4.MN0.G a_n232_43748# 0.0157f
C2620 XA3.XA3.MN0.G a_9848_45156# 6.55e-19
C2621 D<7> a_3440_41284# 6.49e-19
C2622 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MP1.D 0.148f
C2623 XA5.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.D 0.0326f
C2624 XA7.XA6.MP0.G XA7.XA1.XA4.MN0.D 6.07e-19
C2625 XA0.XA9.MN1.G a_920_51492# 6.57e-19
C2626 a_920_52548# XA0.XA7.MP0.G 1.75e-19
C2627 XA7.XA9.MN1.G a_18560_51844# 0.0164f
C2628 a_16040_52196# XA6.XA7.MP0.D 0.0658f
C2629 AVDD a_19928_49732# 0.00159f
C2630 CK_SAMPLE a_5960_50084# 0.00848f
C2631 XA3.XA9.MN1.G XA3.XA8.MP0.D 0.0132f
C2632 a_5960_52196# a_5960_51844# 0.0109f
C2633 a_n232_44452# EN 0.00207f
C2634 a_12368_44452# a_12368_44100# 0.0109f
C2635 XA20.XA2a.MN0.D XA3.XA1.XA4.MP1.D 0.0128f
C2636 XA3.XA1.XA5.MN2.D XA3.XA1.XA2.MP0.D 4.72e-19
C2637 a_11000_51492# XA4.XA6.MP0.G 4.06e-20
C2638 XA2.XA1.XA5.MN2.G XA0.XA6.MP0.G 3.47e-19
C2639 D<2> D<1> 6.86f
C2640 XA8.XA1.XA5.MN2.G a_17408_50436# 0.0046f
C2641 XA4.XA9.MN1.G a_9848_49380# 4.23e-20
C2642 a_7328_52196# VREF 0.00396f
C2643 AVDD a_23600_46564# 0.00159f
C2644 XA20.XA10.MN1.D a_22448_47620# 2.14e-19
C2645 a_19928_51140# a_19928_50788# 0.0109f
C2646 a_12368_43396# a_12368_43044# 0.0109f
C2647 XA1.XA6.MP0.G li_14804_10992# 0.00504f
C2648 XA7.XA6.MP0.G XDAC2.XC32a<0>.XRES16.B 0.00136f
C2649 EN a_11000_42340# 0.159f
C2650 XA7.XA6.MP0.G a_18560_49380# 0.0547f
C2651 XA2.XA1.XA5.MN2.G a_920_47268# 7.1e-20
C2652 XA0.XA7.MP0.G a_2288_47268# 7.1e-20
C2653 AVDD XA6.XA1.XA5.MP0.D 0.159f
C2654 a_22448_50084# a_22448_49732# 0.0109f
C2655 a_8480_49732# a_9848_49732# 8.89e-19
C2656 XA3.XA6.MP0.G a_8480_49028# 0.0137f
C2657 XA20.XA1.MN0.D a_23600_41636# 0.056f
C2658 a_23600_42340# a_23600_41988# 0.0109f
C2659 D<8> li_14804_16116# 0.00508f
C2660 D<3> a_12368_44804# 2.37e-19
C2661 a_11000_48324# a_11000_47972# 0.0109f
C2662 XA3.XA4.MN0.G XA4.XA4.MN0.G 0.12f
C2663 XA20.XA10.MN1.D a_22448_41988# 1.97e-19
C2664 XA20.XA3.MN0.D a_23600_46564# 0.0289f
C2665 AVDD XA5.XA1.XA1.MP1.D 0.0599f
C2666 VREF XA6.XA3.MN0.G 0.608f
C2667 XA3.XA4.MN0.D XA3.XA3.MN0.G 0.158f
C2668 XA5.XA1.XA5.MN2.G a_11000_44100# 0.00556f
C2669 AVDD XA6.XA10.MP0.G 0.853f
C2670 XA0.XA12.MP0.D a_3440_53252# 0.0758f
C2671 XA5.XA11.MN1.G XA4.XA11.MP0.D 0.00856f
C2672 XA8.XA12.MP0.G a_21080_53604# 0.0893f
C2673 DONE a_19928_52900# 9.67e-20
C2674 a_11000_40932# a_11000_40580# 0.0109f
C2675 XA4.XA1.XA1.MN0.D a_9848_40228# 0.00155f
C2676 XA0.XA11.MN1.G XB1.M1.G 0.216f
C2677 XA8.XA1.XA5.MN2.G a_18560_41988# 0.0673f
C2678 XA0.XA7.MP0.G a_2288_41636# 4.13e-19
C2679 a_12368_46564# a_13520_46564# 0.00133f
C2680 a_n232_46564# a_n232_46212# 0.0109f
C2681 XA3.XA4.MN0.G a_7328_44804# 5.54e-19
C2682 XA3.XA3.MN0.G a_7328_46212# 0.155f
C2683 CK_SAMPLE a_4808_50788# 0.157f
C2684 XA1.XA9.MN1.G XA2.XA9.MN1.G 0.0531f
C2685 AVDD a_19928_50436# 0.00154f
C2686 XB1.M1.G a_11000_1390# 0.0684f
C2687 a_12368_2094# a_12368_1742# 0.0109f
C2688 SAR_IN a_13808_1038# 0.00159f
C2689 XB1.XA0.MP0.D a_8408_1742# 0.135f
C2690 XB2.M1.G XB2.XA3.MN1.D 0.015f
C2691 XA20.XA3a.MN0.D a_8480_42692# 0.01f
C2692 a_19928_45156# a_19928_44804# 0.0109f
C2693 a_5960_44804# a_7328_44804# 8.89e-19
C2694 XA5.XA4.MN0.G XA5.XA1.XA4.MN0.D 0.00331f
C2695 XA1.XA3.MN0.G a_3440_43396# 0.00348f
C2696 XA0.XA1.XA5.MN2.D a_n232_44100# 0.0877f
C2697 a_n232_45508# EN 4.27e-19
C2698 SARN XDAC2.X16ab.XRES1B.B 3.59f
C2699 AVDD a_21080_47620# 0.356f
C2700 XA5.XA9.MN1.G XA5.XA6.MP0.D 0.0618f
C2701 li_9184_24300# li_9184_23688# 0.00271f
C2702 XDAC1.X16ab.XRES2.B XDAC1.X16ab.XRES1A.B 0.0136f
C2703 XDAC1.X16ab.XRES4.B XDAC1.XC128b<2>.XRES4.B 0.00284f
C2704 EN a_18560_43044# 5.26e-19
C2705 XA0.XA4.MN0.D XDAC1.XC0.XRES16.B 8.44e-20
C2706 D<2> XDAC1.XC32a<0>.XRES16.B 0.00136f
C2707 XA0.XA6.MP0.G li_14804_20820# 0.00504f
C2708 XA20.XA2a.MN0.D a_14888_41284# 0.0895f
C2709 SARP a_22448_42692# 6.57e-19
C2710 XA8.XA1.XA5.MP1.D a_21080_43396# 0.00176f
C2711 a_21080_43748# XA8.XA1.XA5.MP0.D 0.00176f
C2712 a_9848_43748# a_9848_43396# 0.0109f
C2713 AVDD a_9848_44100# 0.00125f
C2714 a_22448_50436# a_22448_50084# 0.0109f
C2715 XA8.XA1.XA5.MN2.G a_17408_48676# 0.00363f
C2716 XA0.XA7.MP0.G a_920_48324# 0.00455f
C2717 XA3.XA6.MP0.G a_8480_50084# 6.4e-20
C2718 XA3.XA6.MP0.D a_7328_50084# 0.049f
C2719 a_17408_50788# VREF 0.00345f
C2720 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES4.B 0.428f
C2721 XA1.XA3.MN0.G li_14804_26556# 0.00504f
C2722 a_16040_42692# a_16040_42340# 0.0109f
C2723 XA1.XA1.XA4.MN0.D a_3440_42340# 0.0474f
C2724 a_2288_43044# XA1.XA1.XA1.MN0.S 4.06e-20
C2725 XA6.XA1.XA4.MN0.D XA6.XA1.XA4.MP0.D 0.00918f
C2726 EN a_17408_40580# 0.0731f
C2727 XA2.XA1.XA5.MN2.G a_3440_45156# 1.95e-19
C2728 XA8.XA1.XA5.MN2.G XA6.XA1.XA5.MN2.D 6.95e-19
C2729 XA7.XA1.XA5.MN2.G XA7.XA1.XA5.MN2.D 0.0405f
C2730 AVDD a_21080_41988# 0.386f
C2731 XA2.XA6.MP0.G XA1.XA3.MN0.G 0.0307f
C2732 XA20.XA3.MN6.D a_23600_47268# 5.92e-19
C2733 a_22448_49028# a_22448_48676# 0.0109f
C2734 XA5.XA4.MN0.D a_13520_47972# 0.0788f
C2735 VREF a_19928_47972# 7.39e-19
C2736 a_12368_53956# a_13520_53956# 0.00133f
C2737 a_n232_53956# XA0.XA12.MP0.G 0.0704f
C2738 a_920_53956# XA0.XA12.MP0.D 0.0442f
C2739 AVDD a_18560_53604# 0.00166f
C2740 a_14888_54308# XA6.XA11.MN1.G 2.9e-19
C2741 SARP XDAC1.XC32a<0>.XRES1B.B 3.59f
C2742 XA20.XA3a.MN0.D XA20.XA2a.MN0.D 3.6f
C2743 AVDD XB1.XA3.MN1.D 1.65f
C2744 a_17408_47268# a_17408_46916# 0.0109f
C2745 XA4.XA1.XA5.MN2.G a_8480_42692# 1.95e-19
C2746 VREF a_7328_44452# 0.0182f
C2747 XA2.XA4.MN0.D a_4808_44452# 9.25e-20
C2748 a_12368_52900# XA5.XA10.MP0.G 0.0674f
C2749 a_21080_52900# a_22448_52900# 8.89e-19
C2750 XA5.XA10.MP0.D a_12368_52548# 0.00224f
C2751 AVDD a_14888_51140# 0.00166f
C2752 CK_SAMPLE a_11000_51492# 5.02e-19
C2753 a_8408_3150# a_8408_2798# 0.0109f
C2754 a_13808_3502# a_14960_3502# 0.00133f
C2755 XA3.XA1.XA5.MN2.G a_5960_39876# 0.00285f
C2756 XA6.XA3.MN0.G a_16040_44100# 0.00245f
C2757 SARN a_12368_1038# 0.0415f
C2758 XA20.XA3a.MN0.D XA7.XA1.XA2.MP0.D 0.199f
C2759 XA1.XA4.MN0.G a_2288_43044# 0.0222f
C2760 a_2288_51844# XA2.XA1.XA5.MN2.G 8.87e-19
C2761 XA1.XA8.MP0.D a_2288_51492# 0.00224f
C2762 XA4.XA9.MN1.G XA4.XA6.MP2.D 0.0618f
C2763 XA7.XA11.MN1.G VREF 0.39f
C2764 AVDD a_19928_48676# 0.00129f
C2765 CK_SAMPLE a_4808_49028# 7.31e-19
C2766 XA1.XA7.MP0.D a_2288_51140# 0.00224f
C2767 XA6.XA7.MP0.D XA7.XA1.XA5.MN2.G 0.14f
C2768 XA20.XA3a.MN0.D XA5.XA1.XA1.MN0.D 0.0616f
C2769 XA20.XA2a.MN0.D a_23600_42340# 0.00271f
C2770 EN a_13520_43748# 0.00532f
C2771 XA2.XA1.XA5.MP1.D a_5960_43748# 0.049f
C2772 a_7328_50788# XA3.XA6.MP0.G 1.34e-19
C2773 XA20.XA10.MN1.D a_23600_46564# 0.00517f
C2774 a_8480_50436# a_9848_50436# 8.89e-19
C2775 AVDD XA8.XA1.XA5.MN2.D 2.37f
C2776 XA7.XA1.XA5.MN2.G a_17408_49732# 7.1e-20
C2777 XA8.XA1.XA5.MN2.G a_16040_49732# 7.1e-20
C2778 D<1> XA7.XA6.MP0.G 3.47f
C2779 XA0.XA7.MP0.G XA0.XA4.MN0.D 0.123f
C2780 EN a_920_41284# 0.00564f
C2781 XA0.XA1.XA2.MP0.D a_n232_41636# 0.00316f
C2782 XA4.XA1.XA2.MP0.D a_9848_41988# 0.0568f
C2783 XA8.XA1.XA2.MP0.D a_19928_42340# 0.095f
C2784 XA3.XA1.XA4.MP1.D a_7328_42692# 0.049f
C2785 a_19928_43044# a_19928_42692# 0.0109f
C2786 XA20.XA3.MN6.D a_22448_48324# 0.00961f
C2787 a_14888_49380# a_16040_49380# 0.00133f
C2788 XA4.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C2789 XA0.XA7.MP0.G a_2288_46212# 7.1e-20
C2790 XA2.XA1.XA5.MN2.G a_920_46212# 7.1e-20
C2791 XA0.XA6.MP2.G XA3.XA3.MN0.G 0.347f
C2792 D<7> D<8> 0.0324f
C2793 AVDD a_5960_42692# 0.358f
C2794 VREF a_17408_49028# 0.0647f
C2795 XA20.XA9.MP0.D a_22448_44100# 0.0674f
C2796 AVDD a_4808_54308# 0.00166f
C2797 XA20.XA12.MP0.D XA20.XA11.MP0.D 0.0615f
C2798 a_22448_54660# XA20.XA11.MN0.D 0.0215f
C2799 XA20.XA12.MP0.G DONE 0.188f
C2800 a_5960_41636# a_5960_41284# 0.0109f
C2801 a_17408_41636# XA7.XA1.XA1.MN0.S 0.071f
C2802 XA7.XA1.XA5.MN2.G XA6.XA1.XA2.MP0.D 0.144f
C2803 a_9848_47620# a_11000_47620# 0.00133f
C2804 AVDD a_2288_39876# 0.438f
C2805 XA2.XA4.MN0.D a_4808_45508# 9.25e-20
C2806 VREF a_7328_45508# 0.0556f
C2807 D<5> a_7328_43748# 7.77e-20
C2808 XA20.XA3a.MN0.D a_22448_47620# 0.0441f
C2809 a_23600_47972# a_23600_47620# 0.0109f
C2810 XA2.XA4.MN0.G a_5960_46916# 0.0678f
C2811 XA1.XA11.MP0.D a_2288_52900# 0.00176f
C2812 XA4.XA11.MN1.G a_8480_52548# 9.76e-19
C2813 CK_SAMPLE XA7.XA9.MN1.G 0.135f
C2814 AVDD XA7.XA7.MP0.D 1.19f
C2815 DONE a_21080_52196# 0.00421f
C2816 a_3440_53252# XA1.XA10.MP0.D 0.0676f
C2817 a_4808_40228# a_4808_39876# 0.0109f
C2818 XA3.XA6.MP0.G a_8480_42340# 7.76e-20
C2819 a_4808_45860# a_5960_45860# 0.00133f
C2820 XA3.XA3.MN0.G a_8480_45156# 0.0832f
C2821 D<7> a_2288_41284# 7.77e-20
C2822 XA5.XA1.XA5.MN2.G XA5.XA1.XA1.MP1.D 6.68e-19
C2823 XA7.XA6.MP0.G XA7.XA1.XA4.MP0.D 9.97e-19
C2824 XA5.XA10.MP0.G XA6.XA1.XA5.MN2.G 2.18e-19
C2825 XA0.XA9.MN1.G a_n232_51492# 0.0118f
C2826 XA7.XA9.MN1.G a_17408_51844# 6.57e-19
C2827 AVDD a_18560_49732# 0.00159f
C2828 CK_SAMPLE a_4808_50084# 0.167f
C2829 a_14888_52196# XA6.XA7.MP0.D 0.0678f
C2830 a_11000_334# a_11000_n18# 0.0109f
C2831 CK_SAMPLE_BSSW a_14960_n18# 5e-19
C2832 XA0.XA6.MP2.G XDAC1.XC0.XRES2.B 0.00406f
C2833 XA0.XA4.MN0.D a_920_40228# 9.14e-20
C2834 SARN li_14804_16116# 0.00103f
C2835 XA20.XA2a.MN0.D XA2.XA1.XA4.MP1.D 0.0128f
C2836 XA0.XA7.MP0.G XA0.XA6.MP0.G 0.093f
C2837 XA7.XA1.XA5.MN2.G a_17408_50436# 7.1e-20
C2838 XA8.XA1.XA5.MN2.G a_16040_50436# 7.1e-20
C2839 XA8.XA9.MN1.G XA8.XA4.MN0.D 0.00938f
C2840 a_5960_52196# VREF 0.00396f
C2841 D<2> XA6.XA6.MP2.D 0.0399f
C2842 AVDD a_22448_46564# 0.404f
C2843 D<6> a_5960_50788# 0.161f
C2844 XA2.XA6.MN2.D a_4808_50788# 0.0488f
C2845 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES4.B 0.428f
C2846 XA5.XA1.XA2.MP0.D XA5.XA1.XA4.MN1.D 0.056f
C2847 XA20.XA2a.MN0.D a_4808_40228# 2.1e-19
C2848 XA0.XA4.MN0.D li_9184_20820# 0.00504f
C2849 XA0.XA6.MP0.G XDAC2.XC64a<0>.XRES2.B 2.23e-21
C2850 XA7.XA6.MP0.G a_17408_49380# 0.0781f
C2851 XA0.XA7.MP0.G a_920_47268# 0.00363f
C2852 AVDD XA6.XA1.XA5.MN0.D 0.00889f
C2853 XA8.XA1.XA5.MN2.G a_17408_47620# 0.00363f
C2854 a_17408_50084# VREF 0.00382f
C2855 XA3.XA6.MP0.G a_7328_49028# 0.0307f
C2856 XA20.XA1.MN0.D a_22448_41636# 2.43e-19
C2857 a_9848_41988# a_11000_41988# 0.00133f
C2858 XA20.XA3.MN0.D a_22448_46564# 2.46e-19
C2859 AVDD XA4.XA1.XA1.MP1.D 0.0604f
C2860 VREF XA5.XA3.MN0.G 0.608f
C2861 XA8.XA4.MN0.D a_21080_46916# 0.00245f
C2862 XA2.XA4.MN0.D XA3.XA3.MN0.G 0.11f
C2863 XA3.XA4.MN0.D XA2.XA3.MN0.G 0.0258f
C2864 XA5.XA1.XA5.MN2.G a_9848_44100# 2.31e-19
C2865 XA20.XA3.MN6.D a_23600_46212# 0.154f
C2866 a_7328_53604# a_8480_53604# 0.00133f
C2867 AVDD XA5.XA10.MP0.G 0.853f
C2868 XA0.XA12.MP0.D a_2288_53252# 0.0762f
C2869 XA0.XA12.MP0.G a_920_53252# 0.00276f
C2870 XA8.XA12.MP0.G a_19928_53604# 0.1f
C2871 a_22448_40932# a_23600_40932# 0.00133f
C2872 XA8.XA1.XA1.MN0.S a_21080_39876# 2.54e-19
C2873 SARP li_9184_5676# 0.00228f
C2874 XA0.XA7.MP0.G a_920_41636# 0.0756f
C2875 XA8.XA1.XA5.MN2.G a_17408_41988# 0.0734f
C2876 XA7.XA1.XA5.MN2.G a_18560_41988# 0.0039f
C2877 VREF a_21080_43748# 8.43e-19
C2878 D<2> XA6.XA1.XA4.MP0.D 6.08e-19
C2879 CK_SAMPLE a_3440_50788# 0.157f
C2880 XA5.XA10.MP0.G a_13520_52196# 0.0131f
C2881 a_3440_52548# a_3440_52196# 0.0109f
C2882 AVDD a_18560_50436# 0.00154f
C2883 XA1.XA9.MN1.G XA1.XA9.MN0.D 0.034f
C2884 a_14888_52548# XA6.XA9.MN0.D 0.00176f
C2885 a_16040_52548# XA6.XA9.MN1.G 0.0658f
C2886 XB1.M1.G a_9560_1390# 0.0015f
C2887 XB1.XA4.MP0.D a_8408_1390# 0.00559f
C2888 SAR_IN a_12368_1038# 0.0604f
C2889 XB2.M1.G XB2.XA3.MN0.S 0.00399f
C2890 XA20.XA3a.MN0.D a_7328_42692# 0.00443f
C2891 XA6.XA1.XA5.MN2.D a_16040_44452# 0.158f
C2892 XA4.XA6.MP0.G a_11000_40580# 5.5e-19
C2893 XA2.XA4.MN0.D a_5960_41284# 9.14e-20
C2894 XA0.XA6.MP0.G a_920_40228# 5.5e-19
C2895 XA6.XA1.XA5.MN2.G a_13520_51140# 0.0677f
C2896 a_3440_51140# a_4808_51140# 8.89e-19
C2897 AVDD a_19928_47620# 0.00154f
C2898 a_22448_51492# a_22448_51140# 0.0109f
C2899 XA5.XA9.MN1.G XA5.XA6.MP0.G 0.0725f
C2900 XA2.XA7.MP0.D a_4808_50436# 1.37e-19
C2901 XB2.XA4.MP0.D XDAC2.XC1.XRES8.B 0.0129f
C2902 EN a_17408_43044# 0.141f
C2903 XA20.XA2a.MN0.D a_13520_41284# 0.088f
C2904 AVDD a_8480_44100# 0.00125f
C2905 D<6> a_5960_49028# 0.00884f
C2906 XA7.XA1.XA5.MN2.G a_17408_48676# 7.1e-20
C2907 XA8.XA1.XA5.MN2.G a_16040_48676# 7.1e-20
C2908 XA3.XA6.MP0.G a_7328_50084# 0.159f
C2909 a_16040_50788# VREF 0.00345f
C2910 D<2> a_16040_49380# 0.00891f
C2911 D<8> li_14804_26556# 3.5e-20
C2912 XA1.XA1.XA4.MP0.D a_3440_42340# 2.16e-19
C2913 XA1.XA1.XA4.MN0.D a_2288_42340# 2.16e-19
C2914 EN a_16040_40580# 0.0715f
C2915 XA0.XA7.MP0.G a_3440_45156# 1e-19
C2916 XA2.XA1.XA5.MN2.G a_2288_45156# 0.00486f
C2917 AVDD a_19928_41988# 0.00159f
C2918 XA2.XA6.MP0.G D<8> 0.0801f
C2919 XA5.XA6.MP0.G a_13520_46916# 5e-19
C2920 XA20.XA3.MN6.D a_22448_47268# 0.00966f
C2921 XA20.XA3a.MN0.G a_23600_47268# 0.154f
C2922 SARN a_23600_44100# 0.0017f
C2923 XA1.XA6.MP0.G XA3.XA3.MN0.G 0.214f
C2924 a_8480_48676# a_9848_48676# 8.89e-19
C2925 XA5.XA4.MN0.D a_12368_47972# 0.0546f
C2926 VREF a_18560_47972# 7.39e-19
C2927 XA7.XA1.XA5.MN2.G XA6.XA1.XA5.MN2.D 0.108f
C2928 a_n232_53956# XA0.XA12.MP0.D 0.0224f
C2929 AVDD a_17408_53604# 0.383f
C2930 a_13520_54308# XA6.XA11.MN1.G 6.78e-19
C2931 a_13520_41284# XA5.XA1.XA1.MN0.D 0.00224f
C2932 a_2288_41284# a_2288_40932# 0.0109f
C2933 XA2.XA4.MN0.G a_5960_45860# 2.12e-19
C2934 AVDD XB1.XA3.MN0.S 0.183f
C2935 a_3440_46916# a_4808_46916# 8.89e-19
C2936 XA4.XA1.XA5.MN2.G a_7328_42692# 0.00442f
C2937 XA3.XA1.XA5.MN2.G a_8480_42692# 0.0755f
C2938 XA7.XA6.MP0.G XA7.XA1.XA5.MN1.D 7.41e-19
C2939 VREF a_5960_44452# 0.0182f
C2940 XA20.XA3a.MN0.D a_23600_46564# 0.00313f
C2941 a_2288_52900# a_2288_52548# 0.0109f
C2942 AVDD a_13520_51140# 0.00166f
C2943 CK_SAMPLE a_9848_51492# 6.34e-19
C2944 a_14960_3854# a_14960_3502# 0.0109f
C2945 XA6.XA3.MN0.G a_14888_44100# 0.00441f
C2946 SARN a_11000_1038# 0.00166f
C2947 XA20.XA3a.MN0.D XA6.XA1.XA5.MP0.D 7.08e-19
C2948 a_16040_45508# XA6.XA1.XA5.MN2.D 0.0659f
C2949 a_5960_45508# a_5960_45156# 0.0109f
C2950 XA7.XA4.MN0.G a_18560_43396# 0.0104f
C2951 a_13520_51844# a_13520_51492# 0.0109f
C2952 SARN D<7> 0.027f
C2953 XA4.XA9.MN1.G XA4.XA6.MN2.D 0.126f
C2954 XA5.XA12.MP0.G VREF 0.0123f
C2955 AVDD a_18560_48676# 0.00129f
C2956 CK_SAMPLE a_3440_49028# 7.31e-19
C2957 XDAC1.XC0.XRES16.B XDAC1.XC64b<1>.XRES16.B 0.0114f
C2958 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES8.B 0.0228f
C2959 li_9184_29616# li_9184_29004# 0.00271f
C2960 XA20.XA3a.MN0.D XA5.XA1.XA1.MP1.D 0.0093f
C2961 XA0.XA6.MP2.G li_9184_21432# 3.5e-20
C2962 XA20.XA2a.MN0.D a_22448_42340# 0.0092f
C2963 SARN XDAC2.XC1.XRES1A.B 3.59f
C2964 a_14888_44452# XA6.XA1.XA2.MP0.D 5.16e-20
C2965 a_4808_44100# XA2.XA1.XA2.MP0.D 2.92e-19
C2966 XA2.XA1.XA5.MP1.D a_4808_43748# 2.16e-19
C2967 XA2.XA1.XA5.MN1.D a_5960_43748# 2.16e-19
C2968 EN a_12368_43748# 0.166f
C2969 a_18560_44100# a_18560_43748# 0.0109f
C2970 XA20.XA10.MN1.D a_22448_46564# 2.14e-19
C2971 AVDD XA7.XA1.XA5.MN2.D 2.36f
C2972 D<6> a_5960_50084# 0.0155f
C2973 XA7.XA1.XA5.MN2.G a_16040_49732# 0.00457f
C2974 a_22448_51492# VREF 0.00104f
C2975 a_21080_50788# a_21080_50436# 0.0109f
C2976 XDAC1.XC32a<0>.XRES2.B XDAC1.XC32a<0>.XRES16.B 0.457f
C2977 EN a_n232_41284# 0.00433f
C2978 XA0.XA4.MN0.D XDAC1.XC64a<0>.XRES2.B 2.23e-21
C2979 XA1.XA4.MN0.D li_9184_10992# 0.00504f
C2980 XA7.XA1.XA4.MP1.D XA7.XA1.XA4.MN1.D 0.00918f
C2981 XA20.XA3a.MN0.G a_22448_48324# 0.0268f
C2982 XA3.XA6.MP0.G a_8480_47972# 6.28e-19
C2983 XA3.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.51f
C2984 XA0.XA7.MP0.G a_920_46212# 0.00363f
C2985 XA0.XA6.MP2.G XA2.XA3.MN0.G 0.675f
C2986 AVDD a_4808_42692# 0.00125f
C2987 VREF a_16040_49028# 0.0647f
C2988 XA4.XA4.MN0.D a_11000_49028# 0.154f
C2989 a_2288_49380# a_2288_49028# 0.0109f
C2990 AVDD a_3440_54308# 0.00166f
C2991 XA20.XA12.MP0.D DONE 0.0689f
C2992 a_22448_54660# a_23600_54660# 0.00133f
C2993 XA20.XA12.MP0.G XA20.XA11.MN0.D 0.014f
C2994 SARP XDAC1.X16ab.XRES1B.B 3.59f
C2995 VREF a_5960_45508# 0.0556f
C2996 AVDD a_920_39876# 0.44f
C2997 XA20.XA3.MN6.D XA20.XA2.MN1.D 0.014f
C2998 XA1.XA6.MP0.G a_3440_44452# 7.76e-20
C2999 XA2.XA4.MN0.G a_4808_46916# 0.0869f
C3000 XA6.XA1.XA5.MN2.G XA6.XA1.XA2.MP0.D 0.126f
C3001 AVDD XA6.XA7.MP0.D 1.19f
C3002 XA4.XA11.MN1.G a_7328_52548# 7.25e-20
C3003 DONE a_19928_52196# 7.22e-19
C3004 XA8.XA11.MN1.G XA8.XA10.MP0.G 7.66e-19
C3005 XA6.XA11.MP0.D XA6.XA10.MP0.D 0.00986f
C3006 a_2288_53252# XA1.XA10.MP0.D 0.0677f
C3007 a_13520_53252# a_14888_53252# 8.89e-19
C3008 a_16040_40228# a_17408_40228# 8.89e-19
C3009 XA3.XA3.MN0.G a_7328_45156# 0.0546f
C3010 XA5.XA4.MN0.G XA5.XA1.XA5.MN1.D 0.0242f
C3011 XA3.XA6.MP0.G a_7328_42340# 5.5e-19
C3012 a_17408_46212# a_17408_45860# 0.0109f
C3013 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MP1.D 0.144f
C3014 XA0.XA4.MN0.D XA0.XA1.XA4.MP1.D 9.69e-19
C3015 a_22448_52196# a_23600_52196# 0.00133f
C3016 AVDD a_17408_49732# 0.359f
C3017 CK_SAMPLE a_3440_50084# 0.167f
C3018 a_4808_52196# a_4808_51844# 0.0109f
C3019 a_13808_334# a_14960_334# 0.00133f
C3020 CK_SAMPLE_BSSW a_13808_n18# 0.0169f
C3021 a_11000_44452# a_11000_44100# 0.0109f
C3022 SARP a_23600_44100# 0.154f
C3023 XA0.XA4.MN0.D a_n232_40228# 9.25e-20
C3024 XA20.XA2a.MN0.D XA2.XA1.XA4.MN1.D 0.0128f
C3025 XA2.XA4.MN0.G XA2.XA1.XA1.MN0.S 5.22e-20
C3026 XA7.XA1.XA5.MN2.G a_16040_50436# 0.0046f
C3027 D<2> XA6.XA6.MN2.D 1.59e-19
C3028 AVDD a_21080_46564# 0.356f
C3029 a_18560_51140# a_18560_50788# 0.0109f
C3030 XB2.XA3.MN1.D m3_16544_308# 0.0137f
C3031 a_11000_43396# a_11000_43044# 0.0109f
C3032 XA5.XA1.XA2.MP0.D XA5.XA1.XA4.MP1.D 4.34e-19
C3033 XA20.XA2a.MN0.D a_3440_40228# 2.1e-19
C3034 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES8.B 0.00687f
C3035 AVDD XA6.XA1.XA2.MP0.D 0.263f
C3036 XA8.XA1.XA5.MN2.G a_16040_47620# 7.1e-20
C3037 XA7.XA1.XA5.MN2.G a_17408_47620# 7.1e-20
C3038 a_16040_50084# VREF 0.00382f
C3039 a_21080_50084# a_21080_49732# 0.0109f
C3040 a_7328_49732# a_8480_49732# 0.00133f
C3041 D<0> a_21080_48324# 0.0164f
C3042 SARP a_11000_1038# 0.04f
C3043 a_22448_42340# a_22448_41988# 0.0109f
C3044 D<8> XDAC2.XC128a<1>.XRES1A.B 0.00406f
C3045 a_9848_48324# a_9848_47972# 0.0109f
C3046 XA1.XA6.MP0.G a_3440_45508# 7.76e-20
C3047 XA2.XA4.MN0.G XA3.XA4.MN0.G 0.00869f
C3048 a_21080_48324# XA8.XA4.MN0.G 0.0658f
C3049 D<7> SARP 0.137f
C3050 AVDD XA4.XA1.XA1.MN0.D 0.0357f
C3051 VREF XA4.XA3.MN0.G 0.608f
C3052 XA2.XA4.MN0.D XA2.XA3.MN0.G 0.075f
C3053 XA8.XA4.MN0.D a_19928_46916# 0.00396f
C3054 XA1.XA4.MN0.D XA3.XA3.MN0.G 0.113f
C3055 XA3.XA4.MN0.D XA1.XA3.MN0.G 0.0258f
C3056 XA4.XA1.XA5.MN2.G a_9848_44100# 0.0709f
C3057 XA5.XA6.MP0.G a_13520_45860# 1.38e-19
C3058 XA20.XA3.MN6.D a_22448_46212# 0.164f
C3059 AVDD XA4.XA10.MP0.G 0.853f
C3060 XA0.XA12.MP0.G a_n232_53252# 0.0661f
C3061 XA0.XA12.MP0.D a_920_53252# 0.00648f
C3062 XA4.XA11.MN1.G XA4.XA11.MP0.D 0.0102f
C3063 XA3.XA12.MP0.G XA3.XA11.MP0.D 0.0612f
C3064 XA8.XA11.MN1.G a_21080_53604# 0.0658f
C3065 a_9848_40932# a_9848_40580# 0.0109f
C3066 XA8.XA1.XA1.MP1.D a_21080_40580# 0.00176f
C3067 XA3.XA1.XA1.MN0.D a_8480_40228# 0.00155f
C3068 XA8.XA1.XA1.MN0.S a_19928_39876# 2.54e-19
C3069 XA4.XA6.MP0.G a_11000_43044# 5.5e-19
C3070 XA0.XA7.MP0.G a_n232_41636# 0.128f
C3071 XA0.XA11.MN1.G a_13808_2446# 0.00275f
C3072 D<2> XA6.XA1.XA4.MN0.D 0.00144f
C3073 XA0.XA6.MP0.G XA0.XA1.XA4.MP1.D 0.00121f
C3074 XA20.XA3a.MN0.D XA8.XA1.XA5.MN2.D 0.00726f
C3075 a_11000_46564# a_12368_46564# 8.89e-19
C3076 XA2.XA4.MN0.G a_5960_44804# 5.54e-19
C3077 XA2.XA3.MN0.G a_5960_46212# 0.155f
C3078 D<6> a_5960_42340# 7.76e-20
C3079 CK_SAMPLE a_2288_50788# 0.00142f
C3080 XA5.XA10.MP0.G a_12368_52196# 0.0441f
C3081 AVDD a_17408_50436# 0.416f
C3082 a_14888_52548# XA6.XA9.MN1.G 0.0727f
C3083 XB2.XA4.MP0.D a_14960_1742# 0.015f
C3084 XB1.M1.G a_8408_1390# 5.05e-19
C3085 a_11000_2094# a_11000_1742# 0.0109f
C3086 a_14960_2094# XB2.XA0.MP0.D 0.0658f
C3087 SAR_IN a_11000_1038# 9.86e-20
C3088 a_18560_45156# a_18560_44804# 0.0109f
C3089 a_4808_44804# a_5960_44804# 0.00133f
C3090 XA20.XA2a.MN0.D XA0.XA1.XA2.MP0.D 0.223f
C3091 XA6.XA1.XA5.MN2.D a_14888_44452# 0.153f
C3092 XA4.XA6.MP0.G a_9848_40580# 7.76e-20
C3093 XA2.XA4.MN0.D a_4808_41284# 9.25e-20
C3094 SARN li_14804_26556# 0.00103f
C3095 XA0.XA6.MP0.G a_n232_40228# 7.76e-20
C3096 XA20.XA3a.MN0.D a_5960_42692# 0.00443f
C3097 XA6.XA1.XA5.MN2.G a_12368_51140# 0.0754f
C3098 SARN XA2.XA6.MP0.G 0.0551f
C3099 AVDD a_18560_47620# 0.00125f
C3100 a_2288_52900# VREF 0.00396f
C3101 a_7328_51492# D<5> 2.41e-19
C3102 XB1.XA4.MP0.D XDAC1.XC1.XRES2.B 0.00369f
C3103 XDAC2.X16ab.XRES2.B XDAC2.X16ab.XRES16.B 0.457f
C3104 XDAC2.X16ab.XRES8.B XDAC2.X16ab.XRES1A.B 0.0228f
C3105 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES2.B 0.00405f
C3106 D<2> li_9184_13860# 0.00504f
C3107 EN a_16040_43044# 0.141f
C3108 XA20.XA2a.MN0.D a_12368_41284# 0.0685f
C3109 XA3.XA1.XA5.MP0.D XA3.XA1.XA5.MN0.D 0.00918f
C3110 XA8.XA1.XA5.MN1.D a_19928_43396# 0.00176f
C3111 XA3.XA1.XA2.MP0.D XA4.XA1.XA2.MP0.D 0.00435f
C3112 a_19928_43748# XA8.XA1.XA5.MN0.D 0.00176f
C3113 a_8480_43748# a_8480_43396# 0.0109f
C3114 AVDD a_7328_44100# 0.359f
C3115 a_21080_50436# a_21080_50084# 0.0109f
C3116 D<6> a_4808_49028# 5.7e-19
C3117 XA7.XA1.XA5.MN2.G a_16040_48676# 0.00363f
C3118 D<2> a_14888_49380# 5.91e-19
C3119 XDAC2.XC64a<0>.XRES2.B XDAC2.XC1.XRES2.B 1.67e-19
C3120 li_14804_9156# li_14804_8736# 0.00411f
C3121 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES1A.B 0.00405f
C3122 a_14888_42692# a_14888_42340# 0.0109f
C3123 XA1.XA1.XA4.MP0.D a_2288_42340# 0.049f
C3124 XA6.XA1.XA2.MP0.D a_16040_41284# 1.07e-19
C3125 XA2.XA1.XA5.MN2.G a_920_45156# 7.1e-20
C3126 XA0.XA7.MP0.G a_2288_45156# 7.1e-20
C3127 AVDD a_18560_41988# 0.00125f
C3128 XA5.XA6.MP0.G a_12368_46916# 5.5e-19
C3129 XA20.XA3a.MN0.G a_22448_47268# 0.182f
C3130 XA1.XA6.MP0.G XA2.XA3.MN0.G 5.92f
C3131 a_21080_49028# a_21080_48676# 0.0109f
C3132 VREF a_17408_47972# 0.0175f
C3133 XA6.XA1.XA5.MN2.G XA6.XA1.XA5.MN2.D 0.0398f
C3134 a_11000_53956# a_12368_53956# 8.89e-19
C3135 AVDD a_16040_53604# 0.383f
C3136 a_12368_54308# XA6.XA11.MN1.G 8.3e-19
C3137 XA0.XA1.XA1.MN0.S a_920_40580# 0.0318f
C3138 XA5.XA1.XA1.MP2.D a_12368_40932# 0.00176f
C3139 SARP li_9184_16116# 0.00103f
C3140 XA2.XA4.MN0.G a_4808_45860# 0.0146f
C3141 AVDD a_14960_1742# 0.363f
C3142 a_4808_47268# XA2.XA3.MN0.G 2.69e-19
C3143 a_16040_47268# a_16040_46916# 0.0109f
C3144 XA3.XA1.XA5.MN2.G a_7328_42692# 1.97e-19
C3145 XA7.XA6.MP0.G XA7.XA1.XA5.MP1.D 0.00121f
C3146 XA1.XA4.MN0.D a_3440_44452# 9.24e-20
C3147 VREF a_4808_44452# 7.12e-19
C3148 XA20.XA3a.MN0.D a_22448_46564# 0.00881f
C3149 a_11000_52900# XA4.XA10.MP0.G 0.0658f
C3150 a_19928_52900# a_21080_52900# 0.00133f
C3151 XA4.XA10.MP0.D a_11000_52548# 0.00224f
C3152 AVDD a_12368_51140# 0.383f
C3153 CK_SAMPLE a_8480_51492# 6.45e-19
C3154 a_8480_53252# XA3.XA9.MN1.G 5.25e-19
C3155 XA2.XA1.XA5.MN2.G a_4808_39876# 0.00169f
C3156 D<1> a_18560_40932# 5.26e-19
C3157 D<5> a_8480_40580# 5.26e-19
C3158 XA5.XA6.MP0.G XA5.XA1.XA1.MN0.S 0.0146f
C3159 XA20.XA3a.MN0.D XA6.XA1.XA5.MN0.D 0.0106f
C3160 a_14888_45508# XA6.XA1.XA5.MN2.D 0.0674f
C3161 XA7.XA4.MN0.G a_17408_43396# 8.07e-19
C3162 XA0.XA4.MN0.G a_920_43044# 0.0222f
C3163 XA8.XA7.MP0.G a_21080_40228# 0.00361f
C3164 a_920_52196# XA0.XA6.MP2.G 7.56e-20
C3165 XA4.XA9.MN1.G D<4> 0.0378f
C3166 XA6.XA11.MN1.G VREF 0.0162f
C3167 AVDD a_17408_48676# 0.356f
C3168 CK_SAMPLE a_2288_49028# 3.27e-19
C3169 XA0.XA7.MP0.D a_920_51140# 0.00224f
C3170 XA5.XA7.MP0.D XA6.XA1.XA5.MN2.G 0.14f
C3171 XA0.XA8.MP0.D a_920_51492# 0.00224f
C3172 a_920_51844# XA0.XA7.MP0.G 8.87e-19
C3173 XA2.XA3.MN0.G a_4808_41636# 0.00335f
C3174 XA20.XA2a.MN0.D a_21080_42340# 0.00734f
C3175 XA2.XA1.XA5.MN1.D a_4808_43748# 0.0494f
C3176 EN a_11000_43748# 0.166f
C3177 XA20.XA3a.MN0.D XA4.XA1.XA1.MP1.D 0.0093f
C3178 a_7328_50436# a_8480_50436# 0.00133f
C3179 AVDD XA6.XA1.XA5.MN2.D 2.36f
C3180 D<6> a_4808_50084# 5.7e-19
C3181 a_21080_51492# VREF 0.00386f
C3182 XA2.XA1.XA4.MP1.D a_5960_42692# 0.049f
C3183 a_18560_43044# a_18560_42692# 0.0109f
C3184 XA3.XA6.MP0.G a_7328_47972# 8.92e-19
C3185 D<0> a_21080_47268# 0.0148f
C3186 XA6.XA6.MP0.G XA6.XA4.MN0.G 0.0415f
C3187 a_13520_49380# a_14888_49380# 8.89e-19
C3188 XA8.XA1.XA5.MN2.G a_17408_46564# 0.00363f
C3189 XA2.XA1.XA5.MN2.G XA20.XA2a.MN0.D 0.593f
C3190 XA0.XA6.MP2.G XA1.XA3.MN0.G 0.194f
C3191 D<4> a_11000_46916# 0.0185f
C3192 AVDD a_3440_42692# 0.00125f
C3193 XA4.XA4.MN0.D a_9848_49028# 0.156f
C3194 VREF a_14888_49028# 7.81e-19
C3195 AVDD a_2288_54308# 0.448f
C3196 XA20.XA12.MP0.G a_23600_54660# 0.0678f
C3197 XA20.XA12.MP0.D XA20.XA11.MN0.D 0.178f
C3198 a_4808_41636# a_4808_41284# 0.0109f
C3199 a_16040_41636# XA6.XA1.XA1.MP2.D 0.00176f
C3200 XA1.XA1.XA1.MN0.S XA2.XA1.XA1.MN0.S 0.00217f
C3201 XA1.XA4.MN0.D a_3440_45508# 9.24e-20
C3202 XA8.XA4.MN0.D a_19928_45860# 5.88e-20
C3203 AVDD a_n232_39876# 0.00131f
C3204 D<2> XA6.XA1.XA5.MP1.D 7.42e-19
C3205 XA2.XA6.MP0.G SARP 0.0256f
C3206 XA5.XA6.MP0.G a_13520_44804# 7.76e-20
C3207 XA20.XA3a.MN0.G XA20.XA2.MN1.D 0.126f
C3208 XA20.XA3.MN6.D a_23600_45156# 0.134f
C3209 a_22448_47972# a_22448_47620# 0.0109f
C3210 XA1.XA6.MP0.G a_2288_44452# 5.5e-19
C3211 XA8.XA4.MN0.G a_21080_47268# 0.155f
C3212 XA1.XA4.MN0.G a_4808_46916# 2.84e-19
C3213 XA2.XA4.MN0.G a_3440_46916# 2.84e-19
C3214 a_8480_47620# a_9848_47620# 8.89e-19
C3215 XA5.XA1.XA5.MN2.G XA6.XA1.XA2.MP0.D 1.74e-19
C3216 XA6.XA1.XA5.MN2.G XA5.XA1.XA5.MN0.D 7.2e-19
C3217 CK_SAMPLE XA6.XA9.MN1.G 0.134f
C3218 AVDD XA5.XA7.MP0.D 1.19f
C3219 XA0.XA11.MP0.D a_920_52900# 0.00176f
C3220 XA3.XA11.MN1.G a_8480_52548# 0.00103f
C3221 XA8.XA11.MN1.G XA7.XA10.MP0.G 0.00598f
C3222 a_3440_40228# a_3440_39876# 0.0109f
C3223 XA20.XA3a.MN0.D a_8480_44100# 5.04e-20
C3224 XA5.XA4.MN0.G XA5.XA1.XA5.MP1.D 0.00138f
C3225 a_3440_45860# a_4808_45860# 8.89e-19
C3226 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.D 0.0384f
C3227 XA4.XA1.XA5.MN2.G XA4.XA1.XA1.MP1.D 0.00107f
C3228 XA0.XA4.MN0.D XA0.XA1.XA4.MN1.D 9.9e-19
C3229 XA4.XA10.MP0.G XA5.XA1.XA5.MN2.G 2.18e-19
C3230 XA20.XA4.MN0.D a_23600_51492# 0.056f
C3231 AVDD a_16040_49732# 0.359f
C3232 CK_SAMPLE a_2288_50084# 0.00848f
C3233 XA2.XA9.MN1.G XA2.XA8.MP0.D 0.0132f
C3234 a_13520_52196# XA5.XA7.MP0.D 0.0662f
C3235 a_9560_334# a_9560_n18# 0.0109f
C3236 CK_SAMPLE_BSSW a_12368_n18# 7.61e-19
C3237 XA0.XA6.MP2.G li_9184_31872# 0.00508f
C3238 a_22448_44452# a_23600_44452# 0.00133f
C3239 XA20.XA3a.MN0.D a_19928_41988# 0.00547f
C3240 SARN XDAC2.XC128a<1>.XRES1A.B 3.59f
C3241 XA20.XA2a.MN0.D XA1.XA1.XA4.MN1.D 0.0128f
C3242 a_n232_45156# XA0.XA1.XA2.MP0.D 1.56e-20
C3243 XA3.XA9.MN1.G a_8480_49380# 4.23e-20
C3244 D<3> D<1> 0.356f
C3245 AVDD a_19928_46564# 0.00159f
C3246 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC128a<1>.XRES4.B 0.428f
C3247 XB2.XA3.MN1.D m3_16472_308# 0.0137f
C3248 XA6.XA6.MP0.G XDAC2.XC32a<0>.XRES16.B 0.00136f
C3249 XA3.XA3.MN0.G a_9848_39876# 0.0011f
C3250 a_22448_43396# a_23600_43396# 0.00133f
C3251 XA1.XA1.XA2.MP0.D a_3440_42692# 0.0946f
C3252 XA0.XA4.MN0.D XDAC1.XC128b<2>.XRES2.B 0.00405f
C3253 EN a_7328_42340# 0.159f
C3254 XA0.XA6.MP0.G li_14804_10992# 1.85e-20
C3255 XA7.XA1.XA5.MN2.G a_16040_47620# 0.00363f
C3256 AVDD XA5.XA1.XA5.MN0.D 0.00889f
C3257 a_9848_50084# XA4.XA4.MN0.D 3.12e-20
C3258 D<6> a_5960_47972# 0.0147f
C3259 D<3> XA5.XA4.MN0.G 0.26f
C3260 D<0> a_19928_48324# 6.53e-19
C3261 SARP a_9560_1038# 2.97e-20
C3262 a_8480_41988# a_9848_41988# 8.89e-19
C3263 XA1.XA6.MP0.G a_2288_45508# 5.5e-19
C3264 a_19928_48324# XA8.XA4.MN0.G 0.0677f
C3265 XA0.XA6.MP2.G a_920_44452# 1.47e-19
C3266 AVDD XA3.XA1.XA1.MN0.D 0.0357f
C3267 VREF XA3.XA3.MN0.G 0.608f
C3268 XA1.XA4.MN0.D XA2.XA3.MN0.G 0.109f
C3269 XA2.XA4.MN0.D XA1.XA3.MN0.G 0.0258f
C3270 XA3.XA4.MN0.D D<8> 0.0322f
C3271 XA4.XA1.XA5.MN2.G a_8480_44100# 2.31e-19
C3272 XA5.XA6.MP0.G a_12368_45860# 5.5e-19
C3273 XA20.XA3a.MN0.G a_22448_46212# 0.0278f
C3274 a_5960_53604# a_7328_53604# 8.89e-19
C3275 AVDD XA3.XA10.MP0.G 0.853f
C3276 XA0.XA12.MP0.D a_n232_53252# 2.82e-19
C3277 XA4.XA11.MN1.G XA3.XA11.MP0.D 0.0114f
C3278 XA7.XA12.MP0.G a_18560_53604# 0.102f
C3279 XA8.XA11.MN1.G a_19928_53604# 0.0709f
C3280 XA20.XA12.MP0.D a_22448_52900# 1.34e-19
C3281 XA20.XA12.MP0.G a_21080_52900# 7.54e-19
C3282 a_21080_40932# a_22448_40932# 8.89e-19
C3283 XA8.XA1.XA1.MN0.D a_21080_40580# 8.3e-19
C3284 SARP XDAC1.XC1.XRES1A.B 3.59f
C3285 XA4.XA6.MP0.G a_9848_43044# 7.76e-20
C3286 XA0.XA11.MN1.G a_12368_2446# 0.16f
C3287 XA0.XA6.MP0.G XA0.XA1.XA4.MN1.D 7.41e-19
C3288 XA20.XA3a.MN0.D XA7.XA1.XA5.MN2.D 4.79e-19
C3289 XA2.XA4.MN0.G a_4808_44804# 0.00858f
C3290 XA2.XA3.MN0.G a_4808_46212# 0.157f
C3291 D<6> a_4808_42340# 6.49e-19
C3292 XA7.XA1.XA5.MN2.G a_16040_41988# 0.0719f
C3293 CK_SAMPLE a_920_50788# 0.00142f
C3294 a_2288_52548# a_2288_52196# 0.0109f
C3295 AVDD a_16040_50436# 0.416f
C3296 SAR_IP a_12368_1038# 9.86e-20
C3297 a_13808_2094# XB2.XA0.MP0.D 0.0739f
C3298 XA7.XA3.MN0.G XA7.XA1.XA2.MP0.D 0.00212f
C3299 XA20.XA2a.MN0.D a_23600_43748# 0.00246f
C3300 XA20.XA3a.MN0.D a_4808_42692# 0.0099f
C3301 AVDD a_17408_47620# 0.356f
C3302 XA5.XA1.XA5.MN2.G a_12368_51140# 7.1e-20
C3303 XA6.XA1.XA5.MN2.G a_11000_51140# 7.1e-20
C3304 a_2288_51140# a_3440_51140# 0.00133f
C3305 a_21080_51492# a_21080_51140# 0.0109f
C3306 XA8.XA7.MP0.D a_19928_50788# 3.29e-19
C3307 a_920_52900# VREF 0.00396f
C3308 XA1.XA7.MP0.D a_3440_50436# 1.37e-19
C3309 EN a_14888_43044# 6.46e-19
C3310 D<3> XDAC1.XC32a<0>.XRES16.B 0.00136f
C3311 XA20.XA2a.MN0.D a_11000_41284# 0.0669f
C3312 XA3.XA1.XA2.MP0.D XA3.XA1.XA5.MN0.D 0.056f
C3313 a_19928_43748# XA8.XA1.XA2.MP0.D 0.0702f
C3314 D<8> a_n232_40932# 0.00369f
C3315 XA7.XA6.MP0.G XA7.XA6.MP0.D 0.0392f
C3316 AVDD a_5960_44100# 0.359f
C3317 XA2.XA6.MP0.D a_5960_50084# 0.049f
C3318 D<8> XDAC2.XC64b<1>.XRES1A.B 4.06e-21
C3319 a_920_43044# XA0.XA1.XA1.MN0.S 4.06e-20
C3320 XA0.XA7.MP0.G a_920_45156# 0.00486f
C3321 AVDD a_17408_41988# 0.386f
C3322 D<0> a_21080_46212# 0.0202f
C3323 XA1.XA6.MP0.G XA1.XA3.MN0.G 2.44f
C3324 a_7328_48676# a_8480_48676# 0.00133f
C3325 VREF a_16040_47972# 0.0175f
C3326 XA4.XA4.MN0.D a_11000_47972# 0.0546f
C3327 XA0.XA6.MP2.G a_920_45508# 0.00436f
C3328 XA6.XA1.XA5.MN2.G XA5.XA1.XA5.MN2.D 0.108f
C3329 D<4> a_11000_45860# 0.0774f
C3330 CK_SAMPLE a_23600_53956# 0.0683f
C3331 AVDD a_14888_53604# 0.00166f
C3332 a_13520_54308# XA5.XA11.MN1.G 0.00123f
C3333 XA0.XA1.XA1.MN0.S a_n232_40580# 0.00155f
C3334 XA5.XA1.XA1.MN0.S a_12368_40932# 0.0271f
C3335 a_12368_41284# XA5.XA1.XA1.MP1.D 0.00176f
C3336 a_920_41284# a_920_40932# 0.0109f
C3337 XA8.XA4.MN0.G a_21080_46212# 3.46e-19
C3338 XA2.XA4.MN0.G a_3440_45860# 2.2e-19
C3339 XA1.XA4.MN0.G a_4808_45860# 2.2e-19
C3340 XA3.XA6.MP0.G a_8480_43748# 7.76e-20
C3341 AVDD a_13808_1742# 0.00166f
C3342 XA8.XA7.MP0.G XA8.XA1.XA4.MP1.D 0.00353f
C3343 a_2288_46916# a_3440_46916# 0.00133f
C3344 XA3.XA1.XA5.MN2.G a_5960_42692# 0.00442f
C3345 D<1> a_18560_43396# 6.49e-19
C3346 XA1.XA4.MN0.D a_2288_44452# 9.15e-20
C3347 VREF a_3440_44452# 7.12e-19
C3348 D<5> a_8480_43044# 6.49e-19
C3349 XA20.XA3a.MN0.D a_21080_46564# 3.15e-19
C3350 a_920_52900# a_920_52548# 0.0109f
C3351 a_9848_52900# XA4.XA10.MP0.G 0.0681f
C3352 XA4.XA10.MP0.D a_9848_52548# 0.00316f
C3353 AVDD a_11000_51140# 0.383f
C3354 CK_SAMPLE a_7328_51492# 5.02e-19
C3355 XA4.XA11.MN1.G a_8480_51844# 1.13e-19
C3356 DONE XA8.XA7.MP0.G 0.0397f
C3357 a_13808_3854# a_13808_3502# 0.0109f
C3358 XA2.XA1.XA5.MN2.G a_3440_39876# 2.97e-20
C3359 D<5> a_7328_40580# 4.18e-20
C3360 XA5.XA3.MN0.G a_13520_44100# 0.00441f
C3361 XA20.XA3a.MN0.D XA6.XA1.XA2.MP0.D 0.195f
C3362 a_22448_45508# a_23600_45508# 0.00133f
C3363 a_4808_45508# a_4808_45156# 0.0109f
C3364 XA1.XA6.MP0.G a_3440_41284# 3.97e-20
C3365 XA0.XA4.MN0.G a_n232_43044# 0.0409f
C3366 XA8.XA7.MP0.G a_19928_40228# 7.56e-20
C3367 D<1> a_17408_40932# 4.18e-20
C3368 XA4.XA12.MP0.G VREF 0.0119f
C3369 AVDD a_16040_48676# 0.356f
C3370 CK_SAMPLE a_920_49028# 3.27e-19
C3371 XA0.XA7.MP0.D a_n232_51140# 0.00388f
C3372 a_12368_51844# a_12368_51492# 0.0109f
C3373 XA0.XA8.MP0.D a_n232_51492# 0.00224f
C3374 XDAC2.XC64b<1>.XRES1B.B XDAC2.XC64b<1>.XRES4.B 0.428f
C3375 SARN li_14804_6288# 0.00138f
C3376 XA2.XA3.MN0.G a_3440_41636# 4.21e-19
C3377 XA1.XA3.MN0.G a_4808_41636# 4.4e-20
C3378 XA0.XA6.MP2.G XDAC1.XC128b<2>.XRES8.B 4.06e-21
C3379 XA6.XA1.XA5.MN1.D XA6.XA1.XA5.MP1.D 0.00918f
C3380 XA20.XA2a.MN0.D a_19928_42340# 0.0845f
C3381 EN a_9848_43748# 0.00532f
C3382 a_17408_44100# a_17408_43748# 0.0109f
C3383 XA20.XA3a.MN0.D XA4.XA1.XA1.MN0.D 0.0616f
C3384 D<1> XA6.XA6.MP0.G 0.0318f
C3385 AVDD XA5.XA1.XA5.MN2.D 2.36f
C3386 a_19928_50788# a_19928_50436# 0.0109f
C3387 D<2> XA7.XA6.MP0.G 0.112f
C3388 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC64a<0>.XRES1B.B 0.00444f
C3389 li_14804_14472# li_14804_13860# 0.00271f
C3390 XDAC2.XC32a<0>.XRES8.B XDAC2.XC32a<0>.XRES16.B 0.0904f
C3391 XA0.XA4.MN0.D li_9184_10992# 1.85e-20
C3392 XA1.XA4.MN0.D XDAC1.XC64a<0>.XRES8.B 0.00687f
C3393 XA2.XA1.XA4.MP1.D a_4808_42692# 2.16e-19
C3394 XA2.XA1.XA4.MN1.D a_5960_42692# 2.16e-19
C3395 EN XA8.XA1.XA1.MN0.S 0.139f
C3396 D<0> a_19928_47268# 3.18e-19
C3397 XA7.XA1.XA5.MN2.G a_17408_46564# 7.1e-20
C3398 XA8.XA1.XA5.MN2.G a_16040_46564# 7.1e-20
C3399 XA0.XA7.MP0.G XA20.XA2a.MN0.D 0.51f
C3400 XA0.XA6.MP2.G D<8> 1.31f
C3401 D<4> a_9848_46916# 0.00249f
C3402 AVDD a_2288_42692# 0.358f
C3403 a_920_49380# a_920_49028# 0.0109f
C3404 VREF a_13520_49028# 7.81e-19
C3405 AVDD a_920_54308# 0.447f
C3406 a_22448_55012# DONE 1.3e-19
C3407 XA20.XA12.MP0.G a_22448_54660# 0.0739f
C3408 XA20.XA12.MP0.D a_23600_54660# 0.00262f
C3409 a_23600_55012# XA20.XA11.MN0.D 2.39e-19
C3410 a_16040_41636# XA6.XA1.XA1.MN0.S 0.0694f
C3411 XA1.XA1.XA1.MN0.S XA1.XA1.XA1.MP2.D 0.0708f
C3412 SARP li_9184_26556# 0.00103f
C3413 XA1.XA4.MN0.D a_2288_45508# 9.15e-20
C3414 D<2> XA6.XA1.XA5.MN1.D 0.00185f
C3415 AVDD a_23600_40228# 0.00166f
C3416 XA5.XA6.MP0.G a_12368_44804# 5.5e-19
C3417 XA20.XA3a.MN0.G a_23600_45156# 0.0218f
C3418 XA20.XA3.MN6.D a_22448_45156# 0.15f
C3419 XA1.XA4.MN0.G a_3440_46916# 0.0885f
C3420 XA8.XA4.MN0.G a_19928_47268# 0.157f
C3421 XA6.XA1.XA5.MN2.G XA5.XA1.XA5.MP0.D 0.00353f
C3422 AVDD XA4.XA7.MP0.D 1.19f
C3423 XA3.XA11.MN1.G a_7328_52548# 0.00135f
C3424 XA5.XA11.MP0.D XA5.XA10.MP0.D 0.00986f
C3425 a_920_53252# XA0.XA10.MP0.D 0.0661f
C3426 a_12368_53252# a_13520_53252# 0.00133f
C3427 a_14888_40228# a_16040_40228# 0.00133f
C3428 a_16040_46212# a_16040_45860# 0.0109f
C3429 XA8.XA3.MN0.G XA8.XA1.XA5.MN2.D 0.702f
C3430 XA2.XA3.MN0.G a_5960_45156# 0.0546f
C3431 XA4.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.D 0.0288f
C3432 D<4> XA4.XA1.XA1.MN0.S 0.0181f
C3433 XA20.XA9.MP0.D a_23600_51140# 0.00337f
C3434 XA20.XA4.MN0.D a_22448_51492# 2.67e-19
C3435 XA6.XA9.MN0.D a_14888_51844# 0.00176f
C3436 XA6.XA9.MN1.G a_16040_51844# 6.57e-19
C3437 a_21080_52196# a_22448_52196# 8.89e-19
C3438 AVDD a_14888_49732# 0.00159f
C3439 CK_SAMPLE a_920_50084# 0.00848f
C3440 a_3440_52196# a_3440_51844# 0.0109f
C3441 a_12368_52196# XA5.XA7.MP0.D 0.0674f
C3442 a_12368_334# a_13808_334# 8e-19
C3443 CK_SAMPLE_BSSW a_11000_n18# 7.61e-19
C3444 XA20.XA3a.MN0.D a_18560_41988# 0.00547f
C3445 XA20.XA2a.MN0.D XA1.XA1.XA4.MP1.D 0.0128f
C3446 XA2.XA1.XA5.MN2.D XA2.XA1.XA2.MP0.D 4.72e-19
C3447 XA8.XA4.MN0.G a_19928_41636# 6.69e-20
C3448 a_9848_44452# a_9848_44100# 0.0109f
C3449 a_21080_44804# EN 3.4e-19
C3450 SARN XA3.XA4.MN0.D 0.027f
C3451 a_2288_52196# VREF 0.00396f
C3452 AVDD a_18560_46564# 0.00125f
C3453 a_17408_51140# a_17408_50788# 0.0109f
C3454 XA1.XA6.MN2.D a_3440_50788# 0.0488f
C3455 XA3.XA9.MN1.G a_7328_49380# 2.54e-19
C3456 XA7.XA9.MN1.G XA7.XA4.MN0.D 0.00938f
C3457 XA8.XA7.MP0.D a_19928_50084# 7.44e-20
C3458 XB2.XA3.MN1.D m3_26048_1188# 0.17f
C3459 XA3.XA3.MN0.G a_8480_39876# 0.00642f
C3460 a_9848_43396# a_9848_43044# 0.0109f
C3461 XA8.XA1.XA5.MP0.D a_21080_43044# 0.00176f
C3462 XA1.XA1.XA2.MP0.D a_2288_42692# 7.68e-20
C3463 EN a_5960_42340# 0.159f
C3464 XA1.XA6.MP0.G li_14804_11604# 0.00504f
C3465 AVDD XA5.XA1.XA5.MP0.D 0.159f
C3466 a_19928_50084# a_19928_49732# 0.0109f
C3467 a_5960_49732# a_7328_49732# 8.89e-19
C3468 D<6> a_4808_47972# 5.43e-19
C3469 a_21080_42692# XA8.XA1.XA1.MN0.S 6.76e-20
C3470 a_21080_42340# a_21080_41988# 0.0109f
C3471 XA2.XA3.MN0.G XDAC2.XC128a<1>.XRES16.B 3.2e-20
C3472 D<8> li_14804_16728# 0.00508f
C3473 a_8480_48324# a_8480_47972# 0.0109f
C3474 XA1.XA4.MN0.G XA2.XA4.MN0.G 0.12f
C3475 XA0.XA6.MP2.G a_n232_44452# 5.24e-19
C3476 D<4> a_11000_44804# 2.36e-19
C3477 AVDD XA3.XA1.XA1.MP1.D 0.0599f
C3478 VREF XA2.XA3.MN0.G 0.608f
C3479 XA1.XA4.MN0.D XA1.XA3.MN0.G 0.157f
C3480 XA7.XA4.MN0.D a_18560_46916# 0.00396f
C3481 XA0.XA4.MN0.D XA3.XA3.MN0.G 0.123f
C3482 XA2.XA4.MN0.D D<8> 0.0322f
C3483 XA3.XA1.XA5.MN2.G a_8480_44100# 0.0693f
C3484 XA4.XA1.XA5.MN2.G a_7328_44100# 0.00556f
C3485 AVDD XA2.XA10.MP0.G 0.853f
C3486 XA7.XA12.MP0.G a_17408_53604# 0.0877f
C3487 XA8.XA11.MN1.G a_18560_53604# 0.00787f
C3488 a_8480_40932# a_8480_40580# 0.0109f
C3489 XA8.XA1.XA1.MN0.D a_19928_40580# 0.035f
C3490 VREF a_17408_43748# 8.43e-19
C3491 XA0.XA11.MN1.G a_11000_2446# 0.159f
C3492 XA20.XA3a.MN0.D XA6.XA1.XA5.MN2.D 3.88e-19
C3493 a_9848_46564# a_11000_46564# 0.00133f
C3494 XA1.XA4.MN0.G a_4808_44804# 2.2e-19
C3495 XA2.XA4.MN0.G a_3440_44804# 2.2e-19
C3496 XA7.XA1.XA5.MN2.G a_14888_41988# 0.0684f
C3497 CK_SAMPLE a_n232_50788# 0.157f
C3498 AVDD a_14888_50436# 0.00154f
C3499 XA4.XA10.MP0.G a_11000_52196# 0.0441f
C3500 a_13520_52548# XA5.XA9.MN0.D 0.00176f
C3501 XA0.XA9.MN1.G XA1.XA9.MN1.G 0.00217f
C3502 XB1.XA4.MP0.D XB1.XA3.MN1.D 0.376p
C3503 a_14960_2446# XB2.XA3.MN1.D 4.69e-19
C3504 SAR_IP a_11000_1038# 0.0604f
C3505 a_9560_2094# a_9560_1742# 0.0109f
C3506 XB2.M1.G a_14960_1742# 0.0315f
C3507 XB2.XA4.MN0.D a_13808_1742# 0.00176f
C3508 XB2.XA1.MP0.D a_14960_1390# 4.8e-20
C3509 XA5.XA1.XA5.MN2.D a_13520_44452# 0.153f
C3510 D<8> a_n232_43396# 0.00341f
C3511 XA4.XA4.MN0.G XA4.XA1.XA4.MN0.D 0.00331f
C3512 a_17408_45156# a_17408_44804# 0.0109f
C3513 a_3440_44804# a_4808_44804# 8.89e-19
C3514 XA20.XA2a.MN0.D a_22448_43748# 0.00168f
C3515 XA1.XA4.MN0.D a_3440_41284# 9.24e-20
C3516 SARN XDAC2.XC64b<1>.XRES1A.B 3.59f
C3517 XA20.XA3a.MN0.D a_3440_42692# 0.01f
C3518 AVDD a_16040_47620# 0.356f
C3519 XA5.XA1.XA5.MN2.G a_11000_51140# 0.077f
C3520 XA4.XA9.MN1.G XA4.XA6.MP0.D 0.0618f
C3521 XDAC1.X16ab.XRES2.B XDAC1.X16ab.XRES16.B 0.457f
C3522 XDAC1.X16ab.XRES8.B XDAC1.X16ab.XRES1A.B 0.0228f
C3523 XA0.XA6.MP0.G li_14804_21432# 0.00504f
C3524 D<2> XDAC1.XC32a<0>.XRES2.B 0.00405f
C3525 XA20.XA2a.MN0.D a_9848_41284# 0.0895f
C3526 XA3.XA1.XA2.MP0.D XA3.XA1.XA5.MP0.D 4.34e-19
C3527 XA7.XA1.XA5.MN1.D a_18560_43396# 0.00176f
C3528 a_7328_43748# a_7328_43396# 0.0109f
C3529 EN a_13520_43044# 5.26e-19
C3530 a_19928_50436# a_19928_50084# 0.0109f
C3531 a_12368_50788# VREF 0.00345f
C3532 AVDD a_4808_44100# 0.00125f
C3533 XDAC1.XC64a<0>.XRES2.B XDAC1.XC1.XRES2.B 1.67e-19
C3534 li_9184_9156# li_9184_8736# 0.00411f
C3535 XA1.XA3.MN0.G li_14804_27168# 0.00504f
C3536 a_13520_42692# a_13520_42340# 0.0109f
C3537 XA0.XA1.XA4.MP0.D a_920_42340# 0.049f
C3538 XA5.XA1.XA4.MP0.D XA5.XA1.XA4.MN0.D 0.00918f
C3539 EN a_12368_40580# 0.0731f
C3540 XA0.XA7.MP0.G a_n232_45156# 1.95e-19
C3541 AVDD a_16040_41988# 0.386f
C3542 XA0.XA6.MP0.G XA3.XA3.MN0.G 0.326f
C3543 D<0> a_19928_46212# 0.0141f
C3544 XA1.XA6.MP0.G D<8> 0.042f
C3545 a_19928_49028# a_19928_48676# 0.0109f
C3546 XA4.XA4.MN0.D a_9848_47972# 0.0788f
C3547 VREF a_14888_47972# 7.39e-19
C3548 XA0.XA6.MP2.G a_n232_45508# 0.0031f
C3549 XA5.XA1.XA5.MN2.G XA5.XA1.XA5.MN2.D 0.0405f
C3550 XA6.XA1.XA5.MN2.G XA4.XA1.XA5.MN2.D 6.95e-19
C3551 D<4> a_9848_45860# 0.0675f
C3552 a_9848_53956# a_11000_53956# 0.00133f
C3553 a_23600_54308# a_23600_53956# 0.0109f
C3554 CK_SAMPLE a_22448_53956# 0.0766f
C3555 AVDD a_13520_53604# 0.00166f
C3556 a_12368_54308# XA5.XA11.MN1.G 8.45e-19
C3557 SARP XDAC1.XC128a<1>.XRES1A.B 3.59f
C3558 XA8.XA4.MN0.G a_19928_46212# 0.0149f
C3559 XA1.XA4.MN0.G a_3440_45860# 0.0146f
C3560 XA3.XA6.MP0.G a_7328_43748# 5.5e-19
C3561 XA8.XA7.MP0.G XA8.XA1.XA4.MN1.D 7.2e-19
C3562 a_3440_47268# XA1.XA3.MN0.G 2.69e-19
C3563 a_14888_47268# a_14888_46916# 0.0109f
C3564 XA3.XA1.XA5.MN2.G a_4808_42692# 1.95e-19
C3565 XA8.XA1.XA5.MN2.G XA8.XA1.XA4.MP1.D 7.44e-19
C3566 D<1> a_17408_43396# 7.77e-20
C3567 XA20.XA10.MN1.D a_23600_40228# 0.0705f
C3568 XA2.XA1.XA5.MN2.G a_5960_42692# 1.97e-19
C3569 VREF a_2288_44452# 0.0182f
C3570 XA3.XA4.MN0.D SARP 0.0406f
C3571 D<5> a_7328_43044# 7.77e-20
C3572 a_18560_52900# a_19928_52900# 8.89e-19
C3573 XA8.XA11.MN1.G XA7.XA7.MP0.D 4.87e-19
C3574 AVDD a_9848_51140# 0.00166f
C3575 CK_SAMPLE a_5960_51492# 5.02e-19
C3576 a_13808_3854# a_14960_3854# 0.00133f
C3577 XA5.XA3.MN0.G a_12368_44100# 0.00245f
C3578 XA0.XA7.MP0.G a_3440_39876# 0.00325f
C3579 XA2.XA1.XA5.MN2.G a_2288_39876# 8.8e-19
C3580 XA20.XA3a.MN0.D XA5.XA1.XA5.MN0.D 0.0107f
C3581 a_13520_45508# XA5.XA1.XA5.MN2.D 0.0658f
C3582 XA1.XA6.MP0.G a_2288_41284# 4.24e-19
C3583 XA6.XA4.MN0.G a_16040_43396# 8.07e-19
C3584 XA8.XA1.XA5.MN2.G a_19928_40228# 0.0709f
C3585 XA5.XA11.MN1.G VREF 0.39f
C3586 SARN XA0.XA6.MP2.G 0.0343f
C3587 AVDD a_14888_48676# 0.00129f
C3588 CK_SAMPLE a_n232_49028# 7.31e-19
C3589 XA4.XA7.MP0.D XA5.XA1.XA5.MN2.G 0.14f
C3590 XA20.XA2a.MN0.D a_18560_42340# 0.0848f
C3591 XA1.XA3.MN0.G a_3440_41636# 0.00333f
C3592 EN a_8480_43748# 0.00532f
C3593 XA1.XA1.XA5.MN1.D a_3440_43748# 0.0494f
C3594 D<5> li_9184_23076# 0.00504f
C3595 XA20.XA3a.MN0.D XA3.XA1.XA1.MN0.D 0.0616f
C3596 AVDD XA4.XA1.XA5.MN2.D 2.36f
C3597 a_5960_50788# XA2.XA6.MP0.G 1.34e-19
C3598 D<2> XA6.XA6.MP0.D 0.0323f
C3599 a_5960_50436# a_7328_50436# 8.89e-19
C3600 XA3.XA1.XA2.MP0.D a_8480_41988# 0.0568f
C3601 XA7.XA1.XA2.MP0.D a_18560_42340# 0.0966f
C3602 XA2.XA1.XA4.MN1.D a_4808_42692# 0.0474f
C3603 a_17408_43044# a_17408_42692# 0.0109f
C3604 a_12368_49380# a_13520_49380# 0.00133f
C3605 XA7.XA1.XA5.MN2.G a_16040_46564# 0.00363f
C3606 AVDD a_920_42692# 0.358f
C3607 VREF a_12368_49028# 0.0647f
C3608 XA3.XA4.MN0.D a_8480_49028# 0.156f
C3609 a_23600_55012# a_23600_54660# 0.0109f
C3610 XA20.XA12.MP0.D a_22448_54660# 0.0318f
C3611 AVDD a_n232_54308# 0.00166f
C3612 a_3440_41636# a_3440_41284# 0.0109f
C3613 a_14888_41636# XA6.XA1.XA1.MN0.S 0.0674f
C3614 VREF a_2288_45508# 0.0556f
C3615 XA7.XA4.MN0.D a_18560_45860# 5.88e-20
C3616 AVDD a_22448_40228# 0.47f
C3617 XA20.XA3a.MN0.G a_22448_45156# 0.0325f
C3618 a_21080_47972# a_21080_47620# 0.0109f
C3619 XA1.XA4.MN0.G a_2288_46916# 0.0662f
C3620 a_7328_47620# a_8480_47620# 0.00133f
C3621 D<6> a_5960_43748# 7.76e-20
C3622 XA6.XA1.XA5.MN2.G XA5.XA1.XA2.MP0.D 0.146f
C3623 AVDD XA3.XA7.MP0.D 1.19f
C3624 XA0.XA11.MN1.G a_n232_52900# 7.39e-19
C3625 XA3.XA11.MN1.G a_5960_52548# 9.29e-19
C3626 XA7.XA11.MN1.G XA7.XA10.MP0.G 0.0119f
C3627 CK_SAMPLE XA5.XA9.MN1.G 0.135f
C3628 a_n232_53252# XA0.XA10.MP0.D 0.0692f
C3629 a_2288_40228# a_2288_39876# 0.0109f
C3630 a_2288_45860# a_3440_45860# 0.00133f
C3631 XA4.XA4.MN0.G XA4.XA1.XA5.MP1.D 0.00138f
C3632 XA2.XA3.MN0.G a_4808_45156# 0.083f
C3633 XA6.XA6.MP0.G XA6.XA1.XA4.MP0.D 9.97e-19
C3634 XA0.XA6.MP2.G a_920_41284# 7.76e-20
C3635 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.D 0.0825f
C3636 XA3.XA10.MP0.G XA4.XA1.XA5.MN2.G 2.18e-19
C3637 XA6.XA9.MN1.G a_14888_51844# 0.0164f
C3638 AVDD a_13520_49732# 0.00159f
C3639 CK_SAMPLE a_n232_50084# 0.167f
C3640 CK_SAMPLE_BSSW a_9560_n18# 0.0169f
C3641 a_8408_334# a_8408_n18# 0.0109f
C3642 a_21080_44452# a_22448_44452# 8.89e-19
C3643 SARN li_14804_16728# 0.00103f
C3644 XA20.XA2a.MN0.D XA0.XA1.XA4.MP1.D 0.0128f
C3645 XA1.XA4.MN0.G XA1.XA1.XA1.MN0.S 5.22e-20
C3646 a_19928_44804# EN 7.78e-19
C3647 XA0.XA6.MP2.G XDAC1.XC0.XRES8.B 0.00688f
C3648 SARN XA2.XA4.MN0.D 0.027f
C3649 a_920_52196# VREF 0.00396f
C3650 AVDD a_17408_46564# 0.356f
C3651 li_14804_19596# li_14804_19176# 0.00411f
C3652 XDAC2.XC128b<2>.XRES2.B XDAC2.XC128a<1>.XRES2.B 1.67e-19
C3653 XB2.XA3.MN1.D m3_25976_1188# 0.0634f
C3654 XA20.XA2a.MN0.D a_n232_40228# 2.1e-19
C3655 XA0.XA4.MN0.D li_9184_21432# 0.00504f
C3656 a_21080_43396# a_22448_43396# 8.89e-19
C3657 XA0.XA6.MP0.G XDAC2.XC64a<0>.XRES8.B 2.23e-21
C3658 XA6.XA6.MP0.G li_14804_13860# 0.00504f
C3659 AVDD XA5.XA1.XA2.MP0.D 0.263f
C3660 XA2.XA6.MP0.G a_5960_49028# 0.0307f
C3661 a_8480_50084# XA3.XA4.MN0.D 3.12e-20
C3662 a_12368_50084# VREF 0.00382f
C3663 XA6.XA6.MP0.G a_16040_49380# 0.0781f
C3664 a_7328_41988# a_8480_41988# 0.00133f
C3665 D<0> a_21080_45156# 5.9e-19
C3666 a_18560_48324# XA7.XA4.MN0.G 0.0661f
C3667 XA0.XA6.MP2.G SARP 0.312f
C3668 D<4> a_9848_44804# 5.24e-19
C3669 AVDD XA2.XA1.XA1.MP1.D 0.0604f
C3670 VREF XA1.XA3.MN0.G 0.608f
C3671 XA7.XA4.MN0.D a_17408_46916# 0.00245f
C3672 XA0.XA4.MN0.D XA2.XA3.MN0.G 0.11f
C3673 XA1.XA4.MN0.D D<8> 0.0322f
C3674 XA3.XA1.XA5.MN2.G a_7328_44100# 7.1e-20
C3675 XA4.XA1.XA5.MN2.G a_5960_44100# 7.1e-20
C3676 a_4808_53604# a_5960_53604# 0.00133f
C3677 AVDD XA1.XA10.MP0.G 0.853f
C3678 CK_SAMPLE a_23600_53252# 8.74e-19
C3679 XA3.XA11.MN1.G XA3.XA11.MP0.D 0.0383f
C3680 XA2.XA12.MP0.G XA2.XA11.MP0.D 0.0612f
C3681 XA8.XA11.MN1.G a_17408_53604# 0.00979f
C3682 a_19928_40932# a_21080_40932# 0.00133f
C3683 XA7.XA1.XA1.MN0.S a_18560_39876# 2.54e-19
C3684 SARP li_9184_6288# 0.00138f
C3685 VREF a_16040_43748# 8.43e-19
C3686 XA0.XA11.MN1.G a_9560_2446# 0.00275f
C3687 XA20.XA3a.MN0.D XA5.XA1.XA5.MN2.D 4.79e-19
C3688 XA1.XA4.MN0.G a_3440_44804# 0.00858f
C3689 XA8.XA4.MN0.G a_21080_45156# 5.54e-19
C3690 XA1.XA3.MN0.G a_3440_46212# 0.157f
C3691 XA8.XA3.MN0.G a_21080_46564# 0.155f
C3692 XA6.XA1.XA5.MN2.G a_14888_41988# 0.00407f
C3693 AVDD a_13520_50436# 0.00154f
C3694 XA4.XA10.MP0.G a_9848_52196# 0.0131f
C3695 a_920_52548# a_920_52196# 0.0109f
C3696 a_13520_52548# XA5.XA9.MN1.G 0.0711f
C3697 XA0.XA9.MN1.G XA0.XA9.MN0.D 0.034f
C3698 CK_SAMPLE XA8.XA6.MP2.D 0.0158f
C3699 XB1.XA4.MP0.D XB1.XA3.MN0.S 1.67e-19
C3700 XB1.M1.G XB1.XA3.MN1.D 0.015f
C3701 SAR_IP a_9560_1038# 0.00159f
C3702 SAR_IN a_14960_1390# 0.00155f
C3703 XB2.M1.G a_13808_1742# 0.00285f
C3704 a_13808_2094# a_14960_2094# 0.00133f
C3705 XB2.XA1.MP0.D a_13808_1390# 5.87e-20
C3706 XA5.XA1.XA5.MN2.D a_12368_44452# 0.158f
C3707 XA1.XA4.MN0.D a_2288_41284# 9.15e-20
C3708 XA20.XA3a.MN0.D a_2288_42692# 0.00443f
C3709 XA4.XA9.MN1.G XA4.XA6.MN0.D 0.0615f
C3710 a_19928_51492# a_19928_51140# 0.0109f
C3711 AVDD a_14888_47620# 0.00125f
C3712 XA5.XA1.XA5.MN2.G a_9848_51140# 0.0661f
C3713 a_920_51140# a_2288_51140# 8.89e-19
C3714 XA7.XA7.MP0.D a_18560_50788# 3.29e-19
C3715 SARN XA1.XA6.MP0.G 0.171f
C3716 XA20.XA9.MP0.D VREF 0.0259f
C3717 XB2.XA4.MP0.D XDAC2.XC1.XRES4.B 0.00738f
C3718 D<1> XDAC1.XC32a<0>.XRES8.B 4.63e-20
C3719 XA20.XA2a.MN0.D a_8480_41284# 0.088f
C3720 a_18560_43748# XA7.XA1.XA5.MN0.D 0.00176f
C3721 EN a_12368_43044# 0.141f
C3722 XA2.XA6.MN0.D a_4808_50084# 0.0488f
C3723 XA2.XA6.MP0.G a_5960_50084# 0.159f
C3724 a_11000_50788# VREF 0.00345f
C3725 AVDD a_3440_44100# 0.00125f
C3726 D<8> li_14804_27168# 3.5e-20
C3727 XA0.XA1.XA4.MN0.D a_920_42340# 2.16e-19
C3728 XA0.XA1.XA4.MP0.D a_n232_42340# 2.16e-19
C3729 EN a_11000_40580# 0.0715f
C3730 XA2.XA3.MN0.G XDAC2.XC64b<1>.XRES16.B 3.2e-20
C3731 AVDD a_14888_41988# 0.00125f
C3732 XA0.XA6.MP0.G XA2.XA3.MN0.G 0.133f
C3733 a_5960_48676# a_7328_48676# 8.89e-19
C3734 VREF a_13520_47972# 7.39e-19
C3735 XA5.XA1.XA5.MN2.G XA4.XA1.XA5.MN2.D 0.108f
C3736 D<4> a_8480_45860# 1.06e-19
C3737 a_11000_54308# XA5.XA11.MN1.G 0.00177f
C3738 AVDD a_12368_53604# 0.383f
C3739 XA20.XA1.MN0.D a_23600_39876# 1.49e-19
C3740 XA4.XA1.XA1.MP2.D a_11000_40932# 0.00176f
C3741 a_11000_41284# XA4.XA1.XA1.MP1.D 0.00176f
C3742 a_n232_41284# a_n232_40932# 0.0109f
C3743 XA8.XA4.MN0.G a_18560_46212# 2.2e-19
C3744 XA7.XA4.MN0.G a_19928_46212# 2.2e-19
C3745 XA1.XA4.MN0.G a_2288_45860# 2.12e-19
C3746 a_920_46916# a_2288_46916# 8.89e-19
C3747 XA8.XA1.XA5.MN2.G XA8.XA1.XA4.MN1.D 0.0131f
C3748 XA20.XA10.MN1.D a_22448_40228# 0.0658f
C3749 XA2.XA1.XA5.MN2.G a_4808_42692# 0.0739f
C3750 VREF a_920_44452# 0.0182f
C3751 XA2.XA4.MN0.D SARP 0.0536f
C3752 a_n232_52900# a_n232_52548# 0.0109f
C3753 a_8480_52900# XA3.XA10.MP0.G 0.0665f
C3754 XA3.XA10.MP0.D a_8480_52548# 0.00316f
C3755 AVDD a_8480_51140# 0.00166f
C3756 CK_SAMPLE a_4808_51492# 6.34e-19
C3757 XA3.XA11.MN1.G a_8480_51844# 3.12e-19
C3758 XA3.XA4.MN0.D a_8480_42340# 9.24e-20
C3759 SARN a_13808_1390# 9.75e-19
C3760 XA0.XA7.MP0.G a_2288_39876# 0.00278f
C3761 XA20.XA3a.MN0.D XA5.XA1.XA5.MP0.D 7.25e-19
C3762 a_21080_45508# a_22448_45508# 8.89e-19
C3763 a_12368_45508# XA5.XA1.XA5.MN2.D 0.0675f
C3764 a_3440_45508# a_3440_45156# 0.0109f
C3765 XA6.XA4.MN0.G a_14888_43396# 0.0104f
C3766 XA8.XA1.XA5.MN2.G a_18560_40228# 1.34e-19
C3767 XA7.XA1.XA5.MN2.G a_19928_40228# 4.72e-19
C3768 XA3.XA12.MP0.G VREF 0.0123f
C3769 SARN a_23600_51140# 0.16f
C3770 XA3.XA9.MN1.G XA3.XA6.MN2.D 0.126f
C3771 AVDD a_13520_48676# 0.00129f
C3772 a_11000_51844# a_11000_51492# 0.0109f
C3773 XDAC1.XC64b<1>.XRES1B.B XDAC1.XC64b<1>.XRES4.B 0.428f
C3774 a_13520_44452# XA5.XA1.XA2.MP0.D 5.16e-20
C3775 XA20.XA2a.MN0.D a_17408_42340# 0.00768f
C3776 SARN XDAC2.XC1.XRES16.B 55.3f
C3777 XA0.XA6.MP2.G li_9184_22044# 3.5e-20
C3778 a_3440_44100# XA1.XA1.XA2.MP0.D 2.92e-19
C3779 XA1.XA1.XA5.MN1.D a_2288_43748# 2.16e-19
C3780 XA1.XA1.XA5.MP1.D a_3440_43748# 2.16e-19
C3781 EN a_7328_43748# 0.166f
C3782 a_16040_44100# a_16040_43748# 0.0109f
C3783 XA20.XA3a.MN0.D XA3.XA1.XA1.MP1.D 0.0093f
C3784 AVDD XA3.XA1.XA5.MN2.D 2.36f
C3785 XA6.XA1.XA5.MN2.G a_12368_49732# 0.00457f
C3786 D<2> XA6.XA6.MN0.D 0.00148f
C3787 a_17408_51492# VREF 0.00396f
C3788 a_18560_50788# a_18560_50436# 0.0109f
C3789 a_4808_50788# XA2.XA6.MP0.G 1.75e-20
C3790 XDAC1.XC32a<0>.XRES8.B XDAC1.XC32a<0>.XRES16.B 0.0904f
C3791 li_9184_14472# li_9184_13860# 0.00271f
C3792 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC64a<0>.XRES1B.B 0.00444f
C3793 XA0.XA4.MN0.D XDAC1.XC64a<0>.XRES8.B 2.23e-21
C3794 XA7.XA1.XA2.MP0.D a_17408_42340# 2.54e-19
C3795 XA6.XA1.XA4.MN1.D XA6.XA1.XA4.MP1.D 0.00918f
C3796 XA3.XA1.XA2.MP0.D a_7328_41988# 0.0219f
C3797 XA1.XA4.MN0.D li_9184_11604# 0.00504f
C3798 EN XA7.XA1.XA1.MN0.S 0.139f
C3799 XA8.XA6.MP0.G a_21080_48324# 0.00362f
C3800 AVDD a_n232_42692# 0.00125f
C3801 VREF a_11000_49028# 0.0647f
C3802 XA3.XA4.MN0.D a_7328_49028# 0.154f
C3803 a_n232_49380# a_n232_49028# 0.0109f
C3804 a_22448_55364# DONE 5e-20
C3805 XA20.XA12.MP0.D XA20.XA12.MP0.G 0.125f
C3806 AVDD XA20.XA11.MP0.D 0.158f
C3807 SARP XDAC1.XC64b<1>.XRES1A.B 3.59f
C3808 VREF a_920_45508# 0.0556f
C3809 AVDD a_21080_40228# 0.469f
C3810 XA1.XA6.MP0.G SARP 0.026f
C3811 XA7.XA4.MN0.G a_18560_47268# 0.157f
C3812 D<6> a_4808_43748# 6.49e-19
C3813 XA5.XA1.XA5.MN2.G XA5.XA1.XA2.MP0.D 0.126f
C3814 AVDD XA2.XA7.MP0.D 1.19f
C3815 a_4808_53956# XA2.XA9.MN1.G 7.37e-20
C3816 XA7.XA11.MN1.G XA6.XA10.MP0.G 0.0024f
C3817 XA4.XA11.MP0.D XA4.XA10.MP0.D 0.00986f
C3818 a_11000_53252# a_12368_53252# 8.89e-19
C3819 a_13520_40228# a_14888_40228# 8.89e-19
C3820 a_14888_46212# a_14888_45860# 0.0109f
C3821 XA2.XA3.MN0.G a_3440_45156# 2.51e-19
C3822 XA1.XA3.MN0.G a_4808_45156# 4.4e-20
C3823 XA7.XA3.MN0.G XA7.XA1.XA5.MN2.D 0.702f
C3824 XA4.XA4.MN0.G XA4.XA1.XA5.MN1.D 0.0242f
C3825 XA6.XA6.MP0.G XA6.XA1.XA4.MN0.D 6.07e-19
C3826 XA0.XA6.MP2.G a_n232_41284# 6.49e-19
C3827 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MP1.D 0.148f
C3828 XA3.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.D 0.0326f
C3829 XA2.XA6.MP0.G a_5960_42340# 5.5e-19
C3830 XA1.XA9.MN1.G XA1.XA8.MP0.D 0.0132f
C3831 XA6.XA9.MN1.G a_13520_51844# 2.2e-19
C3832 a_19928_52196# a_21080_52196# 0.00133f
C3833 AVDD a_12368_49732# 0.359f
C3834 a_2288_52196# a_2288_51844# 0.0109f
C3835 a_11000_52196# XA4.XA7.MP0.D 0.0658f
C3836 a_11000_334# a_12368_334# 8.89e-19
C3837 CK_SAMPLE_BSSW a_8408_n18# 5e-19
C3838 XA20.XA2a.MN0.D XA0.XA1.XA4.MN1.D 0.0128f
C3839 XA7.XA4.MN0.G a_18560_41636# 6.69e-20
C3840 XA3.XA3.MN0.G a_9848_42692# 7.98e-19
C3841 a_8480_44452# a_8480_44100# 0.0109f
C3842 a_18560_44804# EN 7.78e-19
C3843 XA6.XA1.XA5.MN2.G a_12368_50436# 0.0046f
C3844 SARN XA1.XA4.MN0.D 0.027f
C3845 a_7328_51492# XA3.XA6.MP0.G 4.06e-20
C3846 AVDD a_16040_46564# 0.356f
C3847 a_16040_51140# a_16040_50788# 0.0109f
C3848 XA1.XA6.MP2.D a_2288_50788# 0.049f
C3849 D<3> D<2> 6.37f
C3850 D<4> D<1> 0.0391f
C3851 XA7.XA7.MP0.D a_18560_50084# 7.44e-20
C3852 XB2.XA3.MN1.D m3_16544_1364# 0.0137f
C3853 a_8480_43396# a_8480_43044# 0.0109f
C3854 XA8.XA1.XA5.MN0.D a_19928_43044# 0.00176f
C3855 XA4.XA1.XA2.MP0.D XA4.XA1.XA4.MP1.D 4.34e-19
C3856 XA8.XA1.XA2.MP0.D a_21080_43044# 3.59e-19
C3857 XA5.XA6.MP0.G XDAC2.XC32a<0>.XRES16.B 0.00136f
C3858 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES4.B 0.00405f
C3859 AVDD XA4.XA1.XA5.MP0.D 0.159f
C3860 XA2.XA6.MP0.G a_4808_49028# 0.0137f
C3861 a_11000_50084# VREF 0.00382f
C3862 a_18560_50084# a_18560_49732# 0.0109f
C3863 a_4808_49732# a_5960_49732# 0.00133f
C3864 XA6.XA6.MP0.G a_14888_49380# 0.0547f
C3865 a_19928_42340# a_19928_41988# 0.0109f
C3866 D<8> XDAC2.XC128a<1>.XRES16.B 0.0333f
C3867 D<0> a_19928_45156# 1.28e-19
C3868 a_7328_48324# a_7328_47972# 0.0109f
C3869 XA0.XA4.MN0.G XA1.XA4.MN0.G 0.00869f
C3870 a_17408_48324# XA7.XA4.MN0.G 0.0674f
C3871 AVDD XA2.XA1.XA1.MN0.D 0.0357f
C3872 VREF D<8> 0.608f
C3873 XA0.XA4.MN0.D XA1.XA3.MN0.G 0.11f
C3874 XA3.XA1.XA5.MN2.G a_5960_44100# 0.00556f
C3875 XA7.XA11.MN1.G a_18560_53604# 0.0726f
C3876 AVDD XA0.XA10.MP0.G 0.853f
C3877 CK_SAMPLE a_22448_53252# 0.00809f
C3878 XA3.XA11.MN1.G XA2.XA11.MP0.D 0.00856f
C3879 XA8.XA11.MN1.G a_16040_53604# 9.49e-20
C3880 a_7328_40932# a_7328_40580# 0.0109f
C3881 XA7.XA1.XA1.MN0.D a_18560_40580# 0.035f
C3882 XA7.XA1.XA1.MN0.S a_17408_39876# 2.54e-19
C3883 XA20.XA3a.MN0.D XA4.XA1.XA5.MN2.D 3.88e-19
C3884 a_8480_46564# a_9848_46564# 8.89e-19
C3885 D<3> XA5.XA1.XA4.MN0.D 0.00144f
C3886 XA8.XA4.MN0.G a_19928_45156# 0.00865f
C3887 XA1.XA4.MN0.G a_2288_44804# 5.54e-19
C3888 XA1.XA3.MN0.G a_2288_46212# 0.155f
C3889 XA8.XA3.MN0.G a_19928_46564# 0.156f
C3890 XA6.XA1.XA5.MN2.G a_13520_41988# 0.0673f
C3891 AVDD a_12368_50436# 0.416f
C3892 a_12368_52548# XA5.XA9.MN1.G 0.0674f
C3893 CK_SAMPLE XA8.XA6.MN2.D 0.0548f
C3894 a_8408_2094# a_8408_1742# 0.0109f
C3895 SAR_IN a_13808_1390# 0.00815f
C3896 XB2.M1.G a_12368_1742# 0.00202f
C3897 XB1.M1.G XB1.XA3.MN0.S 0.00399f
C3898 a_13808_2446# XB2.XA3.MN0.S 1.03e-19
C3899 a_16040_45156# a_16040_44804# 0.0109f
C3900 a_2288_44804# a_3440_44804# 0.00133f
C3901 XA20.XA2a.MN0.D a_19928_43748# 4.48e-20
C3902 XA3.XA4.MN0.G XA3.XA1.XA4.MN0.D 0.00331f
C3903 XA3.XA6.MP0.G a_8480_40580# 7.76e-20
C3904 XA7.XA6.MP0.G a_18560_40932# 3.97e-20
C3905 SARN li_14804_27168# 0.00103f
C3906 XA20.XA3a.MN0.D a_920_42692# 0.00443f
C3907 XA4.XA9.MN1.G XA4.XA6.MP0.G 0.0725f
C3908 a_5960_51492# D<6> 2.41e-19
C3909 AVDD a_13520_47620# 0.00125f
C3910 XA8.XA10.MP0.D VREF 0.0119f
C3911 XB1.XA4.MP0.D XDAC1.XC1.XRES8.B 0.0129f
C3912 XDAC2.X16ab.XRES1B.B XDAC2.XC128b<2>.XRES1B.B 0.00444f
C3913 li_14804_24912# li_14804_24300# 0.00271f
C3914 XDAC2.X16ab.XRES8.B XDAC2.X16ab.XRES16.B 0.0904f
C3915 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES1A.B 0.0197f
C3916 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES8.B 0.00687f
C3917 XA20.XA2a.MN0.D a_7328_41284# 0.0685f
C3918 XA7.XA1.XA5.MP1.D a_17408_43396# 0.00176f
C3919 a_5960_43748# a_5960_43396# 0.0109f
C3920 D<4> XDAC1.XC32a<0>.XRES16.B 0.00136f
C3921 EN a_11000_43044# 0.141f
C3922 XA2.XA6.MP0.G a_4808_50084# 6.4e-20
C3923 a_18560_50436# a_18560_50084# 0.0109f
C3924 D<3> a_13520_49380# 5.91e-19
C3925 D<7> a_3440_49028# 5.7e-19
C3926 XA6.XA1.XA5.MN2.G a_12368_48676# 0.00363f
C3927 AVDD a_2288_44100# 0.359f
C3928 XDAC2.XC64a<0>.XRES1A.B XDAC2.XC1.XRES1B.B 0.617f
C3929 a_12368_42692# a_12368_42340# 0.0109f
C3930 XA0.XA1.XA4.MN0.D a_n232_42340# 0.0474f
C3931 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES16.B 0.0282f
C3932 AVDD a_13520_41988# 0.00125f
C3933 XA4.XA6.MP0.G a_11000_46916# 5.5e-19
C3934 XA0.XA6.MP0.G XA1.XA3.MN0.G 2.53f
C3935 XA8.XA6.MP0.G a_21080_47268# 4.52e-20
C3936 a_18560_49028# a_18560_48676# 0.0109f
C3937 VREF a_12368_47972# 0.0175f
C3938 XA3.XA4.MN0.D a_8480_47972# 0.0788f
C3939 XA4.XA1.XA5.MN2.G XA4.XA1.XA5.MN2.D 0.0398f
C3940 AVDD a_11000_53604# 0.383f
C3941 DONE XA20.XA10.MN0.D 7.2e-19
C3942 a_8480_53956# a_9848_53956# 8.89e-19
C3943 a_22448_54308# a_22448_53956# 0.0109f
C3944 a_9848_54308# XA5.XA11.MN1.G 2.54e-19
C3945 XA20.XA1.MN0.D a_22448_39876# 2.54e-19
C3946 XA4.XA1.XA1.MN0.S a_11000_40932# 0.0271f
C3947 a_22448_41284# a_23600_41284# 0.00133f
C3948 SARP li_9184_16728# 0.00103f
C3949 AVDD a_9560_1742# 0.00166f
C3950 XA7.XA4.MN0.G a_18560_46212# 0.0149f
C3951 XA6.XA6.MP0.G XA6.XA1.XA5.MP1.D 0.00121f
C3952 a_13520_47268# a_13520_46916# 0.0109f
C3953 XA8.XA1.XA5.MN2.G XA7.XA1.XA4.MN1.D 7.2e-19
C3954 XA2.XA1.XA5.MN2.G a_3440_42692# 1.95e-19
C3955 XA0.XA4.MN0.D a_920_44452# 9.14e-20
C3956 XA1.XA4.MN0.D SARP 0.169f
C3957 VREF a_n232_44452# 7.12e-19
C3958 XA7.XA11.MN1.G XA7.XA7.MP0.D 0.00283f
C3959 a_7328_52900# XA3.XA10.MP0.G 0.0674f
C3960 a_17408_52900# a_18560_52900# 0.00133f
C3961 XA3.XA10.MP0.D a_7328_52548# 0.00224f
C3962 AVDD a_7328_51140# 0.383f
C3963 CK_SAMPLE a_3440_51492# 6.45e-19
C3964 XA3.XA11.MN1.G a_7328_51844# 4.48e-19
C3965 XA4.XA3.MN0.G a_11000_44100# 0.00245f
C3966 XA3.XA4.MN0.D a_7328_42340# 9.15e-20
C3967 SARN a_12368_1390# 0.0415f
C3968 XA20.XA3a.MN0.D XA5.XA1.XA2.MP0.D 0.199f
C3969 XA7.XA1.XA5.MN2.G a_18560_40228# 0.0825f
C3970 XA8.XA1.XA5.MN2.G a_17408_40228# 0.00255f
C3971 XA0.XA7.MP0.G a_920_39876# 0.00285f
C3972 XA4.XA11.MN1.G VREF 0.0162f
C3973 XA3.XA9.MN1.G XA3.XA6.MP2.D 0.0618f
C3974 AVDD a_12368_48676# 0.356f
C3975 CK_SAMPLE a_22448_49380# 2.27e-19
C3976 XA3.XA7.MP0.D XA4.XA1.XA5.MN2.G 0.14f
C3977 XA20.XA2a.MN0.D a_16040_42340# 0.00732f
C3978 XA1.XA1.XA5.MP1.D a_2288_43748# 0.049f
C3979 EN a_5960_43748# 0.166f
C3980 D<5> XDAC1.X16ab.XRES1A.B 0.00405f
C3981 XA20.XA3a.MN0.D XA2.XA1.XA1.MP1.D 0.0093f
C3982 AVDD XA2.XA1.XA5.MN2.D 2.36f
C3983 D<3> XA7.XA6.MP0.G 0.123f
C3984 XA6.XA1.XA5.MN2.G a_11000_49732# 7.1e-20
C3985 XA5.XA1.XA5.MN2.G a_12368_49732# 7.1e-20
C3986 D<7> a_3440_50084# 5.7e-19
C3987 D<2> XA6.XA6.MP0.G 2.21f
C3988 a_16040_51492# VREF 0.00396f
C3989 D<1> XA5.XA6.MP0.G 0.0318f
C3990 a_4808_50436# a_5960_50436# 0.00133f
C3991 XA1.XA1.XA4.MN1.D a_3440_42692# 0.0474f
C3992 a_16040_43044# a_16040_42692# 0.0109f
C3993 a_11000_49380# a_12368_49380# 8.89e-19
C3994 AVDD XA8.XA1.XA4.MP1.D 0.0991f
C3995 XA2.XA6.MP0.G a_5960_47972# 8.92e-19
C3996 VREF a_9848_49028# 7.81e-19
C3997 XA5.XA6.MP0.G XA5.XA4.MN0.G 0.0415f
C3998 XA8.XA6.MP0.G a_19928_48324# 0.00245f
C3999 a_22448_55012# a_22448_54660# 0.0109f
C4000 a_23600_55012# XA20.XA12.MP0.G 0.0658f
C4001 AVDD DONE 2.49f
C4002 a_2288_41636# a_2288_41284# 0.0109f
C4003 XA0.XA1.XA1.MN0.S XA1.XA1.XA1.MN0.S 0.00217f
C4004 AVDD a_19928_40228# 0.00166f
C4005 XA0.XA4.MN0.D a_920_45508# 9.14e-20
C4006 XA0.XA6.MP0.G a_920_44452# 5.5e-19
C4007 a_19928_47972# a_19928_47620# 0.0109f
C4008 XA0.XA4.MN0.G a_920_46916# 0.0678f
C4009 XA7.XA4.MN0.G a_17408_47268# 0.155f
C4010 a_5960_47620# a_7328_47620# 8.89e-19
C4011 XA5.XA1.XA5.MN2.G XA4.XA1.XA5.MP0.D 0.00353f
C4012 AVDD XA1.XA7.MP0.D 1.19f
C4013 a_23600_53604# XA20.XA9.MP0.D 4.23e-19
C4014 CK_SAMPLE XA4.XA9.MN1.G 0.134f
C4015 a_920_40228# a_920_39876# 0.0109f
C4016 a_920_45860# a_2288_45860# 8.89e-19
C4017 XA20.XA3a.MN0.D a_3440_44100# 5.04e-20
C4018 XA1.XA3.MN0.G a_3440_45156# 0.0832f
C4019 XA3.XA1.XA5.MN2.G XA3.XA1.XA1.MP1.D 6.68e-19
C4020 XA2.XA6.MP0.G a_4808_42340# 7.76e-20
C4021 XA5.XA9.MN1.G a_14888_51844# 2.2e-19
C4022 XA5.XA9.MN0.D a_13520_51844# 0.00176f
C4023 XA2.XA10.MP0.G XA3.XA1.XA5.MN2.G 2.18e-19
C4024 XA8.XA10.MP0.G a_19928_51492# 6.8e-20
C4025 AVDD a_11000_49732# 0.359f
C4026 a_9848_52196# XA4.XA7.MP0.D 0.0678f
C4027 CK_SAMPLE XA20.XA3.MN6.D 8.52e-20
C4028 CK_SAMPLE_BSSW a_14960_334# 0.0679f
C4029 a_19928_44452# a_21080_44452# 0.00133f
C4030 XA20.XA3a.MN0.D a_14888_41988# 0.00547f
C4031 SARN XDAC2.XC128a<1>.XRES16.B 55.3f
C4032 XA20.XA2a.MN0.D a_23600_43044# 0.00257f
C4033 XA8.XA1.XA5.MN2.D a_21080_43748# 0.00388f
C4034 XA3.XA3.MN0.G a_8480_42692# 0.00343f
C4035 a_17408_44804# EN 3.4e-19
C4036 XA0.XA6.MP2.G li_9184_32484# 0.00508f
C4037 D<3> XA5.XA6.MN2.D 1.59e-19
C4038 XA5.XA1.XA5.MN2.G a_12368_50436# 7.1e-20
C4039 XA6.XA1.XA5.MN2.G a_11000_50436# 7.1e-20
C4040 AVDD a_14888_46564# 0.00125f
C4041 D<7> a_2288_50788# 0.161f
C4042 XA2.XA9.MN1.G a_5960_49380# 2.54e-19
C4043 XA6.XA9.MN1.G XA6.XA4.MN0.D 0.00938f
C4044 li_9184_19596# li_9184_19176# 0.00411f
C4045 XDAC1.XC128b<2>.XRES2.B XDAC1.XC128a<1>.XRES2.B 1.67e-19
C4046 XB2.XA3.MN1.D m3_16472_1364# 0.0137f
C4047 a_19928_43396# a_21080_43396# 0.00133f
C4048 XA8.XA1.XA2.MP0.D a_19928_43044# 0.0292f
C4049 XA4.XA1.XA2.MP0.D XA4.XA1.XA4.MN1.D 0.056f
C4050 XA0.XA4.MN0.D XDAC1.XC128b<2>.XRES8.B 0.00687f
C4051 EN a_2288_42340# 0.159f
C4052 XA0.XA6.MP0.G li_14804_11604# 1.85e-20
C4053 XA6.XA6.MP0.G XDAC2.XC32a<0>.XRES2.B 0.00405f
C4054 AVDD XA4.XA1.XA5.MN0.D 0.00889f
C4055 D<1> a_18560_48324# 6.53e-19
C4056 XA6.XA1.XA5.MN2.G a_12368_47620# 0.00363f
C4057 D<4> XA4.XA4.MN0.G 0.26f
C4058 SARP a_12368_1390# 0.00463f
C4059 a_5960_41988# a_7328_41988# 8.89e-19
C4060 XA4.XA6.MP0.G a_11000_45860# 5.5e-19
C4061 AVDD XA1.XA1.XA1.MN0.D 0.0357f
C4062 XA0.XA4.MN0.D D<8> 0.0813f
C4063 XA6.XA4.MN0.D a_16040_46916# 0.00245f
C4064 XA8.XA7.MP0.G a_22448_44452# 0.00104f
C4065 XA3.XA1.XA5.MN2.G a_4808_44100# 2.31e-19
C4066 XA0.XA6.MP0.G a_920_45508# 5.5e-19
C4067 XA7.XA11.MN1.G a_17408_53604# 0.073f
C4068 XA6.XA12.MP0.G a_16040_53604# 0.0893f
C4069 AVDD a_23600_52900# 0.0232f
C4070 CK_SAMPLE a_21080_53252# 6.94e-19
C4071 a_3440_53604# a_4808_53604# 8.89e-19
C4072 a_18560_40932# a_19928_40932# 8.89e-19
C4073 XA7.XA1.XA1.MN0.D a_17408_40580# 8.3e-19
C4074 SARP XDAC1.XC1.XRES16.B 55.3f
C4075 XA7.XA6.MP0.G a_18560_43396# 7.76e-20
C4076 XA20.XA3a.MN0.D XA3.XA1.XA5.MN2.D 4.79e-19
C4077 D<3> XA5.XA1.XA4.MP0.D 6.09e-19
C4078 XA0.XA11.MN1.G XB2.XA1.MP0.D 0.0452f
C4079 XA3.XA6.MP0.G a_8480_43044# 7.76e-20
C4080 XA7.XA4.MN0.G a_19928_45156# 2.2e-19
C4081 XA8.XA4.MN0.G a_18560_45156# 2.2e-19
C4082 XA3.XA3.MN0.G XA20.XA2a.MN0.D 0.271f
C4083 D<7> a_3440_42340# 6.49e-19
C4084 XA5.XA1.XA5.MN2.G a_13520_41988# 0.0039f
C4085 XA6.XA1.XA5.MN2.G a_12368_41988# 0.0734f
C4086 AVDD a_11000_50436# 0.416f
C4087 XA3.XA10.MP0.G a_8480_52196# 0.0131f
C4088 a_n232_52548# a_n232_52196# 0.0109f
C4089 CK_SAMPLE D<0> 0.0537f
C4090 XB2.XA1.MN0.D a_13808_1390# 3.62e-20
C4091 SAR_IN a_12368_1390# 0.0597f
C4092 a_12368_2094# a_13808_2094# 8e-19
C4093 a_9560_2094# XB1.XA0.MP0.D 0.0723f
C4094 XA20.XA2a.MN0.D a_18560_43748# 2.91e-20
C4095 XA4.XA1.XA5.MN2.D a_11000_44452# 0.158f
C4096 XA6.XA3.MN0.G XA6.XA1.XA2.MP0.D 0.00212f
C4097 XA3.XA6.MP0.G a_7328_40580# 5.5e-19
C4098 XA7.XA6.MP0.G a_17408_40932# 4.24e-19
C4099 XA20.XA3a.MN0.D a_n232_42692# 0.00984f
C4100 XA0.XA7.MP0.D a_n232_50436# 1.37e-19
C4101 a_18560_51492# a_18560_51140# 0.0109f
C4102 AVDD a_12368_47620# 0.356f
C4103 XA4.XA1.XA5.MN2.G a_8480_51140# 0.0677f
C4104 a_n232_51140# a_920_51140# 0.00133f
C4105 XA20.XA9.MP0.D a_23600_49732# 0.00334f
C4106 XA7.XA10.MP0.D VREF 0.0118f
C4107 XA20.XA2a.MN0.D a_5960_41284# 0.0669f
C4108 a_18560_43748# XA7.XA1.XA2.MP0.D 0.0686f
C4109 a_17408_43748# XA7.XA1.XA5.MP0.D 0.00176f
C4110 D<6> XDAC1.XC32a<0>.XRES1A.A 0.0138f
C4111 EN a_9848_43044# 6.46e-19
C4112 D<3> a_12368_49380# 0.00891f
C4113 D<7> a_2288_49028# 0.00884f
C4114 XA5.XA1.XA5.MN2.G a_12368_48676# 7.1e-20
C4115 XA6.XA1.XA5.MN2.G a_11000_48676# 7.1e-20
C4116 XA6.XA6.MP0.G XA7.XA6.MP0.G 7.36f
C4117 AVDD a_920_44100# 0.359f
C4118 D<8> XDAC2.XC64b<1>.XRES16.B 3.84e-19
C4119 AVDD a_12368_41988# 0.386f
C4120 D<5> a_9848_45860# 1.06e-19
C4121 XA4.XA6.MP0.G a_9848_46916# 5e-19
C4122 XA0.XA6.MP0.G D<8> 5.44f
C4123 a_4808_48676# a_5960_48676# 0.00133f
C4124 VREF a_11000_47972# 0.0175f
C4125 XA3.XA4.MN0.D a_7328_47972# 0.0546f
C4126 XA8.XA7.MP0.G a_22448_45508# 6.64e-19
C4127 XA4.XA1.XA5.MN2.G XA3.XA1.XA5.MN2.D 0.108f
C4128 AVDD a_9848_53604# 0.00166f
C4129 DONE XA20.XA10.MN1.D 0.0422f
C4130 XA20.XA11.MN0.D XA20.XA10.MN0.D 0.0708f
C4131 XA8.XA1.XA1.MP2.D XA8.XA1.XA1.MP1.D 0.0488f
C4132 a_9848_41284# XA4.XA1.XA1.MN0.D 0.00224f
C4133 XA7.XA4.MN0.G a_17408_46212# 3.46e-19
C4134 XA0.XA4.MN0.G a_920_45860# 2.12e-19
C4135 XA6.XA6.MP0.G XA6.XA1.XA5.MN1.D 7.41e-19
C4136 a_n232_46916# a_920_46916# 0.00133f
C4137 XA7.XA1.XA5.MN2.G XA7.XA1.XA4.MN1.D 0.0131f
C4138 XA8.XA1.XA5.MN2.G XA7.XA1.XA4.MP1.D 0.00353f
C4139 XA2.XA1.XA5.MN2.G a_2288_42692# 0.00442f
C4140 XA0.XA7.MP0.G a_3440_42692# 0.0755f
C4141 XA0.XA4.MN0.D a_n232_44452# 9.25e-20
C4142 AVDD a_8408_1742# 0.363f
C4143 XA20.XA9.MP0.D XA20.XA4.MN0.D 0.037f
C4144 AVDD a_5960_51140# 0.383f
C4145 CK_SAMPLE a_2288_51492# 5.02e-19
C4146 a_4808_53252# XA2.XA9.MN1.G 5.25e-19
C4147 XA3.XA11.MN1.G a_5960_51844# 2.62e-19
C4148 XA0.XA11.MN1.G SARN 0.393f
C4149 XA7.XA11.MN1.G XA6.XA7.MP0.D 8.25e-19
C4150 XA4.XA3.MN0.G a_9848_44100# 0.00441f
C4151 SARN a_11000_1390# 0.012f
C4152 D<2> a_16040_40932# 4.07e-20
C4153 XA20.XA3a.MN0.D XA4.XA1.XA5.MP0.D 7.08e-19
C4154 a_19928_45508# a_21080_45508# 0.00133f
C4155 a_11000_45508# XA4.XA1.XA5.MN2.D 0.0659f
C4156 a_2288_45508# a_2288_45156# 0.0109f
C4157 XA5.XA4.MN0.G a_13520_43396# 0.0104f
C4158 D<6> a_5960_40580# 4.07e-20
C4159 XA7.XA1.XA5.MN2.G a_17408_40228# 0.0128f
C4160 XA4.XA6.MP0.G XA4.XA1.XA1.MN0.S 0.0172f
C4161 XA20.XA9.MP0.D a_23600_50436# 0.00643f
C4162 XA2.XA12.MP0.G VREF 0.0119f
C4163 XA3.XA9.MN1.G D<5> 0.0378f
C4164 AVDD a_11000_48676# 0.356f
C4165 CK_SAMPLE a_21080_49380# 2.21e-19
C4166 a_9848_51844# a_9848_51492# 0.0109f
C4167 XA8.XA7.MP0.D a_21080_51492# 0.0893f
C4168 XDAC2.XC0.XRES2.B XDAC2.XC64b<1>.XRES2.B 1.67e-19
C4169 li_14804_30036# li_14804_29616# 0.00411f
C4170 XA0.XA6.MP2.G XDAC1.XC128b<2>.XRES4.B 4.06e-21
C4171 XA5.XA1.XA5.MP1.D XA5.XA1.XA5.MN1.D 0.00918f
C4172 XA20.XA2.MN1.D a_23600_43396# 0.0604f
C4173 XA20.XA2a.MN0.D a_14888_42340# 0.0843f
C4174 SARN li_14804_6900# 0.00117f
C4175 EN a_4808_43748# 0.00532f
C4176 a_14888_44100# a_14888_43748# 0.0109f
C4177 XA20.XA3a.MN0.D XA2.XA1.XA1.MN0.D 0.0616f
C4178 AVDD XA1.XA1.XA5.MN2.D 2.36f
C4179 XA5.XA1.XA5.MN2.G a_11000_49732# 0.00457f
C4180 D<7> a_2288_50084# 0.0155f
C4181 a_17408_50788# a_17408_50436# 0.0109f
C4182 XDAC2.XC32a<0>.XRES8.B XDAC2.XC32a<0>.XRES2.B 0.44f
C4183 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES16.B 0.0483f
C4184 XA1.XA1.XA4.MN1.D a_2288_42692# 2.16e-19
C4185 XA1.XA1.XA4.MP1.D a_3440_42692# 2.16e-19
C4186 XA1.XA4.MN0.D XDAC1.XC64a<0>.XRES4.B 0.00405f
C4187 XA0.XA4.MN0.D li_9184_11604# 1.85e-20
C4188 EN XA6.XA1.XA1.MN0.S 0.139f
C4189 D<1> a_18560_47268# 3.18e-19
C4190 AVDD XA8.XA1.XA4.MN1.D 0.00926f
C4191 XA2.XA6.MP0.G a_4808_47972# 6.28e-19
C4192 XA2.XA4.MN0.D a_5960_49028# 0.154f
C4193 VREF a_8480_49028# 7.81e-19
C4194 D<5> a_8480_46916# 0.00249f
C4195 a_22448_55012# XA20.XA12.MP0.G 0.0725f
C4196 a_23600_55012# XA20.XA12.MP0.D 0.0215f
C4197 AVDD XA20.XA11.MN0.D 0.679f
C4198 a_12368_41636# XA5.XA1.XA1.MP2.D 0.00176f
C4199 a_13520_41636# XA5.XA1.XA1.MN0.S 0.0658f
C4200 XA0.XA1.XA1.MN0.S XA0.XA1.XA1.MP2.D 0.0708f
C4201 SARP li_9184_27168# 0.00103f
C4202 AVDD a_18560_40228# 0.00131f
C4203 XA0.XA6.MP0.G a_n232_44452# 7.76e-20
C4204 D<3> XA5.XA1.XA5.MN1.D 0.00185f
C4205 XA0.XA4.MN0.G a_n232_46916# 0.0869f
C4206 XA5.XA1.XA5.MN2.G XA4.XA1.XA5.MN0.D 7.2e-19
C4207 XA4.XA6.MP0.G a_11000_44804# 5.5e-19
C4208 XA0.XA4.MN0.D a_n232_45508# 9.25e-20
C4209 XA2.XA11.MN1.G a_4808_52548# 2.85e-19
C4210 XA6.XA11.MN1.G XA6.XA10.MP0.G 7.66e-19
C4211 XA20.XA10.MN1.D a_23600_52900# 0.0779f
C4212 XA3.XA11.MP0.D XA3.XA10.MP0.D 0.00986f
C4213 a_9848_53252# a_11000_53252# 0.00133f
C4214 AVDD XA0.XA7.MP0.D 1.19f
C4215 a_12368_40228# a_13520_40228# 0.00133f
C4216 a_13520_46212# a_13520_45860# 0.0109f
C4217 XA6.XA3.MN0.G XA6.XA1.XA5.MN2.D 0.702f
C4218 XA1.XA3.MN0.G a_2288_45156# 0.0546f
C4219 XA3.XA4.MN0.G XA3.XA1.XA5.MN1.D 0.0242f
C4220 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MP1.D 0.144f
C4221 D<1> a_18560_41636# 6.49e-19
C4222 XA5.XA9.MN1.G a_13520_51844# 0.0164f
C4223 a_18560_52196# a_19928_52196# 8.89e-19
C4224 AVDD a_9848_49732# 0.00159f
C4225 a_920_52196# a_920_51844# 0.0109f
C4226 CK_SAMPLE XA20.XA3a.MN0.G 0.00455f
C4227 a_9560_334# a_11000_334# 8e-19
C4228 CK_SAMPLE_BSSW a_13808_334# 0.0816f
C4229 a_14960_686# a_14960_334# 0.0109f
C4230 XA20.XA3a.MN0.D a_13520_41988# 0.00547f
C4231 XA1.XA1.XA5.MN2.D XA1.XA1.XA2.MP0.D 4.72e-19
C4232 XA20.XA2a.MN0.D a_22448_43044# 0.00366f
C4233 XA8.XA1.XA5.MN2.D a_19928_43748# 0.00224f
C4234 XA0.XA4.MN0.G XA0.XA1.XA1.MN0.S 5.22e-20
C4235 a_7328_44452# a_7328_44100# 0.0109f
C4236 a_16040_44804# EN 3.4e-19
C4237 D<3> XA5.XA6.MP2.D 0.0399f
C4238 XA5.XA1.XA5.MN2.G a_11000_50436# 0.0046f
C4239 SARN XA0.XA4.MN0.D 0.027f
C4240 XA20.XA9.MP0.D a_23600_48676# 0.00334f
C4241 AVDD a_13520_46564# 0.00125f
C4242 a_14888_51140# a_14888_50788# 0.0109f
C4243 XA2.XA9.MN1.G a_4808_49380# 4.23e-20
C4244 XB2.XA3.MN1.D m3_26048_2244# 0.17f
C4245 a_7328_43396# a_7328_43044# 0.0109f
C4246 XA0.XA1.XA2.MP0.D a_920_42692# 7.68e-20
C4247 XA7.XA6.MP0.G XDAC2.XC32a<0>.XRES8.B 4.63e-20
C4248 XA2.XA3.MN0.G a_4808_39876# 0.00627f
C4249 EN a_920_42340# 0.159f
C4250 XA1.XA6.MP0.G li_14804_12216# 0.00504f
C4251 AVDD XA4.XA1.XA2.MP0.D 0.263f
C4252 D<1> a_17408_48324# 0.0164f
C4253 XA6.XA1.XA5.MN2.G a_11000_47620# 7.1e-20
C4254 XA5.XA1.XA5.MN2.G a_12368_47620# 7.1e-20
C4255 XA0.XA11.MN1.G SARP 0.523f
C4256 a_17408_50084# a_17408_49732# 0.0109f
C4257 a_3440_49732# a_4808_49732# 8.89e-19
C4258 D<7> a_3440_47972# 5.43e-19
C4259 SARP a_11000_1390# 0.0396f
C4260 a_18560_42340# a_18560_41988# 0.0109f
C4261 D<8> li_14804_17340# 0.00508f
C4262 a_16040_48324# XA6.XA4.MN0.G 0.0658f
C4263 XA4.XA6.MP0.G a_9848_45860# 1.38e-19
C4264 AVDD XA1.XA1.XA1.MP1.D 0.0599f
C4265 VREF a_22448_46916# 0.001f
C4266 XA6.XA4.MN0.D a_14888_46916# 0.00396f
C4267 XA8.XA7.MP0.G a_21080_44452# 0.00486f
C4268 XA0.XA6.MP0.G a_n232_45508# 7.76e-20
C4269 XA2.XA1.XA5.MN2.G a_4808_44100# 0.0709f
C4270 a_5960_48324# a_5960_47972# 0.0109f
C4271 XA7.XA11.MN1.G a_16040_53604# 0.0124f
C4272 XA6.XA12.MP0.G a_14888_53604# 0.1f
C4273 XA1.XA12.MP0.G XA1.XA11.MP0.D 0.0612f
C4274 AVDD a_22448_52900# 0.486f
C4275 XA2.XA11.MN1.G XA2.XA11.MP0.D 0.0102f
C4276 a_5960_40932# a_5960_40580# 0.0109f
C4277 XA7.XA1.XA1.MP1.D a_17408_40580# 0.00176f
C4278 XA2.XA1.XA1.MN0.D a_4808_40228# 0.00155f
C4279 VREF a_12368_43748# 8.43e-19
C4280 XA3.XA4.MN0.D a_8480_43748# 9.24e-20
C4281 XA20.XA3a.MN0.D XA2.XA1.XA5.MN2.D 3.88e-19
C4282 a_7328_46564# a_8480_46564# 0.00133f
C4283 XA0.XA11.MN1.G SAR_IN 0.377f
C4284 XA3.XA6.MP0.G a_7328_43044# 5.5e-19
C4285 XA7.XA4.MN0.G a_18560_45156# 0.00865f
C4286 XA0.XA4.MN0.G a_920_44804# 5.54e-19
C4287 XA2.XA3.MN0.G XA20.XA2a.MN0.D 0.26f
C4288 D<8> a_920_46212# 0.155f
C4289 XA7.XA3.MN0.G a_18560_46564# 0.156f
C4290 D<7> a_2288_42340# 7.77e-20
C4291 XA7.XA6.MP0.G a_17408_43396# 5.5e-19
C4292 AVDD a_9848_50436# 0.00154f
C4293 XA3.XA10.MP0.G a_7328_52196# 0.0441f
C4294 CK_SAMPLE XA7.XA6.MN2.D 0.039f
C4295 a_8408_2094# XB1.XA0.MP0.D 0.0674f
C4296 XB2.XA4.MP0.D XB2.XA0.MP0.D 0.134f
C4297 SAR_IN a_11000_1390# 1.31e-19
C4298 a_14888_45156# a_14888_44804# 0.0109f
C4299 a_920_44804# a_2288_44804# 8.89e-19
C4300 XA4.XA1.XA5.MN2.D a_9848_44452# 0.153f
C4301 XA0.XA4.MN0.D a_920_41284# 9.14e-20
C4302 SARN XDAC2.XC64b<1>.XRES16.B 55.3f
C4303 XA20.XA3a.MN0.D XA8.XA1.XA4.MP1.D 3.4e-19
C4304 AVDD a_11000_47620# 0.356f
C4305 XA4.XA1.XA5.MN2.G a_7328_51140# 0.0754f
C4306 XA6.XA10.MP0.D VREF 0.0118f
C4307 SARN XA0.XA6.MP0.G 0.392f
C4308 XDAC1.X16ab.XRES1B.B XDAC1.XC128b<2>.XRES1B.B 0.00444f
C4309 li_9184_24912# li_9184_24300# 0.00271f
C4310 XDAC1.X16ab.XRES8.B XDAC1.X16ab.XRES16.B 0.0904f
C4311 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES1A.B 0.0197f
C4312 XA20.XA2a.MN0.D a_4808_41284# 0.0895f
C4313 XA2.XA1.XA5.MN0.D XA2.XA1.XA5.MP0.D 0.00918f
C4314 XA6.XA1.XA5.MP1.D a_16040_43396# 0.00176f
C4315 a_4808_43748# a_4808_43396# 0.0109f
C4316 D<2> XDAC1.XC32a<0>.XRES8.B 4.63e-20
C4317 EN a_8480_43044# 5.26e-19
C4318 XA0.XA6.MP0.G li_14804_22044# 0.00504f
C4319 a_17408_50436# a_17408_50084# 0.0109f
C4320 XA5.XA1.XA5.MN2.G a_11000_48676# 0.00363f
C4321 XA1.XA6.MN0.D a_3440_50084# 0.0488f
C4322 XA6.XA6.MP0.G XA6.XA6.MP0.D 0.0392f
C4323 a_7328_50788# VREF 0.00345f
C4324 AVDD a_n232_44100# 0.00125f
C4325 XDAC1.XC64a<0>.XRES1A.B XDAC1.XC1.XRES1B.B 0.617f
C4326 a_11000_42692# a_11000_42340# 0.0109f
C4327 a_23600_42692# XA20.XA1.MN0.D 0.00176f
C4328 XA4.XA1.XA4.MN0.D XA4.XA1.XA4.MP0.D 0.00918f
C4329 XA5.XA1.XA2.MP0.D a_12368_41284# 1.07e-19
C4330 EN a_7328_40580# 0.0731f
C4331 XA1.XA3.MN0.G li_14804_27780# 0.00504f
C4332 AVDD a_11000_41988# 0.386f
C4333 D<5> a_8480_45860# 0.0675f
C4334 a_17408_49028# a_17408_48676# 0.0109f
C4335 VREF a_9848_47972# 7.39e-19
C4336 XA8.XA7.MP0.G a_21080_45508# 0.00595f
C4337 XA3.XA1.XA5.MN2.G XA3.XA1.XA5.MN2.D 0.0405f
C4338 XA4.XA1.XA5.MN2.G XA2.XA1.XA5.MN2.D 6.95e-19
C4339 D<1> a_18560_46212# 0.0141f
C4340 AVDD a_8480_53604# 0.00166f
C4341 XA20.XA11.MN0.D XA20.XA10.MN1.D 0.342f
C4342 DONE XA8.XA12.MP0.G 0.00304f
C4343 a_7328_53956# a_8480_53956# 0.00133f
C4344 a_21080_54308# a_21080_53956# 0.0109f
C4345 a_9848_54308# XA4.XA11.MN1.G 2.9e-19
C4346 XA8.XA1.XA1.MN0.S XA8.XA1.XA1.MP1.D 0.0615f
C4347 a_21080_41284# a_22448_41284# 8.89e-19
C4348 SARP XDAC1.XC128a<1>.XRES16.B 55.3f
C4349 XA0.XA4.MN0.G a_n232_45860# 0.0146f
C4350 a_n232_47268# D<8> 2.69e-19
C4351 a_12368_47268# a_12368_46916# 0.0109f
C4352 D<6> a_5960_43044# 7.76e-20
C4353 XA7.XA1.XA5.MN2.G XA7.XA1.XA4.MP1.D 7.44e-19
C4354 XA0.XA7.MP0.G a_2288_42692# 1.97e-19
C4355 XA0.XA4.MN0.D SARP 0.391f
C4356 AVDD XB2.XA0.MP0.D 2.28f
C4357 D<2> a_16040_43396# 7.76e-20
C4358 XA2.XA6.MP0.G a_5960_43748# 5.5e-19
C4359 XA2.XA10.MP0.D a_5960_52548# 0.00224f
C4360 a_16040_52900# a_17408_52900# 8.89e-19
C4361 a_5960_52900# XA2.XA10.MP0.G 0.0658f
C4362 AVDD a_4808_51140# 0.00166f
C4363 CK_SAMPLE a_920_51492# 5.02e-19
C4364 a_8408_3150# a_9560_3150# 0.00133f
C4365 XA3.XA3.MN0.G a_9848_44100# 7.98e-19
C4366 XA2.XA4.MN0.D a_5960_42340# 9.14e-20
C4367 XA0.XA6.MP0.G a_920_41284# 4.24e-19
C4368 D<2> a_14888_40932# 5.24e-19
C4369 XA20.XA3a.MN0.D XA4.XA1.XA5.MN0.D 0.0106f
C4370 a_9848_45508# XA4.XA1.XA5.MN2.D 0.0674f
C4371 XA5.XA4.MN0.G a_12368_43396# 8.07e-19
C4372 D<6> a_4808_40580# 5.24e-19
C4373 XA7.XA1.XA5.MN2.G a_16040_40228# 0.0108f
C4374 XA20.XA9.MP0.D a_22448_50436# 1.26e-19
C4375 XA3.XA11.MN1.G VREF 0.39f
C4376 AVDD a_9848_48676# 0.00129f
C4377 CK_SAMPLE a_19928_49380# 8.18e-19
C4378 XA2.XA7.MP0.D XA3.XA1.XA5.MN2.G 0.14f
C4379 XA8.XA7.MP0.D a_19928_51492# 0.124f
C4380 XA20.XA2.MN1.D a_22448_43396# 0.0553f
C4381 XA20.XA2a.MN0.D a_13520_42340# 0.0848f
C4382 D<8> a_n232_41636# 0.00335f
C4383 EN a_3440_43748# 0.00532f
C4384 XA0.XA1.XA5.MP1.D a_920_43748# 0.049f
C4385 XA20.XA3a.MN0.D XA1.XA1.XA1.MN0.D 0.0616f
C4386 XA20.XA9.MP0.D a_23600_47620# 0.00334f
C4387 AVDD XA0.XA1.XA5.MN2.D 2.36f
C4388 a_3440_50436# a_4808_50436# 8.89e-19
C4389 XA1.XA1.XA4.MP1.D a_2288_42692# 0.049f
C4390 a_14888_43044# a_14888_42692# 0.0109f
C4391 XA6.XA1.XA5.MN2.G a_12368_46564# 0.00363f
C4392 a_9848_49380# a_11000_49380# 0.00133f
C4393 D<1> a_17408_47268# 0.0148f
C4394 AVDD XA7.XA1.XA4.MN1.D 0.00889f
C4395 VREF a_7328_49028# 0.0647f
C4396 XA2.XA4.MN0.D a_4808_49028# 0.156f
C4397 D<5> a_7328_46916# 0.0185f
C4398 a_22448_55012# XA20.XA12.MP0.D 0.0313f
C4399 AVDD a_23600_54660# 0.00159f
C4400 a_920_41636# a_920_41284# 0.0109f
C4401 a_12368_41636# XA5.XA1.XA1.MN0.S 0.071f
C4402 AVDD a_17408_40228# 0.464f
C4403 XA0.XA6.MP0.G SARP 0.0267f
C4404 a_18560_47972# a_18560_47620# 0.0109f
C4405 D<3> XA5.XA1.XA5.MP1.D 7.43e-19
C4406 XA6.XA4.MN0.G a_16040_47268# 0.155f
C4407 a_4808_47620# a_5960_47620# 0.00133f
C4408 XA5.XA1.XA5.MN2.G XA4.XA1.XA2.MP0.D 0.144f
C4409 XA4.XA6.MP0.G a_9848_44804# 7.76e-20
C4410 XA6.XA4.MN0.D a_14888_45860# 5.88e-20
C4411 VREF a_22448_45860# 0.0013f
C4412 XA2.XA11.MN1.G a_3440_52548# 9.76e-19
C4413 CK_SAMPLE XA3.XA9.MN1.G 0.135f
C4414 XA6.XA11.MN1.G XA5.XA10.MP0.G 0.00598f
C4415 XA20.XA10.MN1.D a_22448_52900# 0.0661f
C4416 XA8.XA11.MP0.D a_21080_53252# 0.0494f
C4417 AVDD a_23600_52196# 0.00193f
C4418 a_n232_40228# a_n232_39876# 0.0109f
C4419 a_n232_45860# a_920_45860# 0.00133f
C4420 XA8.XA7.MP0.G a_22448_41284# 9.75e-19
C4421 XA3.XA4.MN0.G XA3.XA1.XA5.MP1.D 0.00138f
C4422 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.D 0.0384f
C4423 D<1> a_17408_41636# 7.77e-20
C4424 XA2.XA1.XA5.MN2.G XA2.XA1.XA1.MP1.D 0.00107f
C4425 D<5> XA3.XA1.XA1.MN0.S 0.0133f
C4426 XA1.XA10.MP0.G XA2.XA1.XA5.MN2.G 2.18e-19
C4427 XA0.XA9.MN1.G XA0.XA8.MP0.D 0.0132f
C4428 XA7.XA10.MP0.G a_18560_51492# 6.8e-20
C4429 AVDD a_8480_49732# 0.00159f
C4430 a_8480_52196# XA3.XA7.MP0.D 0.0662f
C4431 CK_SAMPLE XA8.XA6.MP0.D 0.00103f
C4432 XA5.XA9.MN1.G a_12368_51844# 6.57e-19
C4433 CK_SAMPLE_BSSW a_12368_334# 5.73e-19
C4434 a_18560_44452# a_19928_44452# 8.89e-19
C4435 SARN li_14804_17340# 0.00103f
C4436 XA20.XA2a.MN0.D a_21080_43044# 0.00168f
C4437 a_14888_44804# EN 7.78e-19
C4438 XA0.XA6.MP2.G XDAC1.XC0.XRES4.B 0.00406f
C4439 D<5> D<1> 0.0013f
C4440 D<4> D<2> 0.269f
C4441 SARN a_23600_49732# 0.163f
C4442 XA8.XA9.MN1.G VREF 0.0728f
C4443 XA20.XA9.MP0.D a_22448_48676# 0.073f
C4444 AVDD a_12368_46564# 0.356f
C4445 XA0.XA6.MP2.D a_920_50788# 0.049f
C4446 XDAC2.XC128b<2>.XRES1A.B XDAC2.XC128a<1>.XRES1B.B 0.617f
C4447 XB2.XA3.MN1.D m3_25976_2244# 0.0634f
C4448 a_18560_43396# a_19928_43396# 8.89e-19
C4449 XA7.XA1.XA5.MN0.D a_18560_43044# 0.00176f
C4450 XA0.XA1.XA2.MP0.D a_n232_42692# 0.0962f
C4451 XA20.XA2a.MN0.D a_19928_40580# 0.00138f
C4452 XA0.XA4.MN0.D li_9184_22044# 0.00504f
C4453 XA4.XA6.MP0.G XDAC2.XC32a<0>.XRES16.B 0.00136f
C4454 XA2.XA3.MN0.G a_3440_39876# 4.21e-19
C4455 XA1.XA3.MN0.G a_4808_39876# 4.4e-20
C4456 EN a_n232_42340# 0.00568f
C4457 XA0.XA6.MP0.G XDAC2.XC64a<0>.XRES4.B 2.23e-21
C4458 AVDD XA3.XA1.XA5.MN0.D 0.00889f
C4459 a_4808_50084# XA2.XA4.MN0.D 3.12e-20
C4460 a_7328_50084# VREF 0.00382f
C4461 D<7> a_2288_47972# 0.0147f
C4462 XA5.XA1.XA5.MN2.G a_11000_47620# 0.00363f
C4463 SARP a_9560_1390# 9.75e-19
C4464 a_17408_42692# XA7.XA1.XA1.MN0.S 6.76e-20
C4465 a_4808_41988# a_5960_41988# 0.00133f
C4466 a_14888_48324# XA6.XA4.MN0.G 0.0677f
C4467 AVDD XA0.XA1.XA1.MP1.D 0.0604f
C4468 VREF a_21080_46916# 0.0536f
C4469 XA8.XA7.MP0.G a_19928_44452# 1.86e-19
C4470 D<5> a_8480_44804# 5.26e-19
C4471 XA2.XA1.XA5.MN2.G a_3440_44100# 2.31e-19
C4472 XA2.XA11.MN1.G XA1.XA11.MP0.D 0.0114f
C4473 XA7.XA11.MN1.G a_14888_53604# 0.00305f
C4474 AVDD a_21080_52900# 0.387f
C4475 a_2288_53604# a_3440_53604# 0.00133f
C4476 a_17408_40932# a_18560_40932# 0.00133f
C4477 XA6.XA1.XA1.MN0.S a_16040_39876# 2.54e-19
C4478 SARP li_9184_6900# 0.00117f
C4479 XA20.XA3a.MN0.D XA1.XA1.XA5.MN2.D 4.79e-19
C4480 XA0.XA11.MN1.G XB2.XA1.MN0.D 0.00904f
C4481 XA0.XA4.MN0.G a_n232_44804# 0.00858f
C4482 XA7.XA4.MN0.G a_17408_45156# 5.54e-19
C4483 XA1.XA3.MN0.G XA20.XA2a.MN0.D 0.265f
C4484 D<8> a_n232_46212# 0.157f
C4485 XA7.XA3.MN0.G a_17408_46564# 0.155f
C4486 XA5.XA1.XA5.MN2.G a_11000_41988# 0.0719f
C4487 XA3.XA4.MN0.D a_7328_43748# 9.15e-20
C4488 VREF a_11000_43748# 8.43e-19
C4489 AVDD a_8480_50436# 0.00154f
C4490 DONE a_21080_50788# 4.11e-19
C4491 XA20.XA4.MN0.D SARN 0.304f
C4492 a_9848_52548# XA4.XA9.MN0.D 0.00176f
C4493 a_11000_52548# XA4.XA9.MN1.G 0.0658f
C4494 a_22448_52548# a_23600_52548# 0.00133f
C4495 CK_SAMPLE XA7.XA6.MP2.D 3.06e-19
C4496 SAR_IP a_12368_1390# 1.31e-19
C4497 a_11000_2094# a_12368_2094# 8.89e-19
C4498 XB1.XA4.MN0.D a_9560_1742# 0.00176f
C4499 XB2.XA4.MN0.D XB2.XA0.MP0.D 0.012f
C4500 XA0.XA4.MN0.D a_n232_41284# 9.25e-20
C4501 XA20.XA3a.MN0.D XA8.XA1.XA4.MN1.D 3.4e-19
C4502 XA3.XA1.XA5.MN2.G a_7328_51140# 7.1e-20
C4503 XA4.XA1.XA5.MN2.G a_5960_51140# 7.1e-20
C4504 XA6.XA7.MP0.D a_14888_50788# 3.29e-19
C4505 a_17408_51492# a_17408_51140# 0.0109f
C4506 AVDD a_9848_47620# 0.00125f
C4507 XA5.XA10.MP0.D VREF 0.0118f
C4508 XA3.XA9.MN1.G XA3.XA6.MN0.D 0.0615f
C4509 SARN a_23600_50436# 0.0189f
C4510 XB2.XA4.MP0.D XDAC2.XC1.XRES1B.B 0.00184f
C4511 XA20.XA2a.MN0.D a_3440_41284# 0.088f
C4512 XA2.XA1.XA2.MP0.D XA2.XA1.XA5.MP0.D 4.34e-19
C4513 EN a_7328_43044# 0.141f
C4514 XA20.XA9.MP0.D XA20.XA2a.MN0.D 0.0338f
C4515 D<0> XA8.XA4.MN0.D 0.203f
C4516 a_5960_50788# VREF 0.00345f
C4517 AVDD a_23600_44452# 0.00154f
C4518 EN a_5960_40580# 0.0715f
C4519 D<8> li_14804_27780# 3.5e-20
C4520 XA8.XA4.MN0.D XA8.XA4.MN0.G 0.708f
C4521 AVDD a_9848_41988# 0.00125f
C4522 D<5> a_7328_45860# 0.0774f
C4523 a_3440_48676# a_4808_48676# 8.89e-19
C4524 XA2.XA4.MN0.D a_5960_47972# 0.0546f
C4525 VREF a_8480_47972# 7.39e-19
C4526 XA8.XA7.MP0.G a_19928_45508# 2.31e-19
C4527 XA3.XA1.XA5.MN2.G XA2.XA1.XA5.MN2.D 0.108f
C4528 D<1> a_17408_46212# 0.0202f
C4529 AVDD a_7328_53604# 0.383f
C4530 a_23600_54660# XA20.XA10.MN1.D 4.3e-19
C4531 a_8480_54308# XA4.XA11.MN1.G 6.78e-19
C4532 XA8.XA1.XA1.MN0.S XA8.XA1.XA1.MN0.D 0.0743f
C4533 a_8480_41284# XA3.XA1.XA1.MN0.D 0.00224f
C4534 XA7.XA1.XA5.MN2.G XA6.XA1.XA4.MP1.D 0.00353f
C4535 D<6> a_4808_43044# 6.49e-19
C4536 XA6.XA4.MN0.G a_16040_46212# 3.46e-19
C4537 XA0.XA7.MP0.G a_920_42692# 0.00442f
C4538 VREF a_22448_44804# 0.00165f
C4539 AVDD XB1.XA0.MP0.D 2.28f
C4540 D<2> a_14888_43396# 6.49e-19
C4541 XA2.XA6.MP0.G a_4808_43748# 7.76e-20
C4542 XA20.XA3.MN0.D a_23600_44452# 0.0764f
C4543 XA20.XA10.MN1.D a_23600_52196# 0.00486f
C4544 XA2.XA10.MP0.D a_4808_52548# 0.00316f
C4545 a_4808_52900# XA2.XA10.MP0.G 0.0681f
C4546 XA8.XA10.MP0.D XA8.XA10.MP0.G 0.194f
C4547 AVDD a_3440_51140# 0.00166f
C4548 CK_SAMPLE a_n232_51492# 6.34e-19
C4549 XB1.XA2.MN0.G a_9560_3150# 0.0674f
C4550 XA3.XA3.MN0.G a_8480_44100# 0.00776f
C4551 XA0.XA6.MP0.G a_n232_41284# 3.97e-20
C4552 XA20.XA3a.MN0.D XA4.XA1.XA2.MP0.D 0.195f
C4553 a_18560_45508# a_19928_45508# 8.89e-19
C4554 a_920_45508# a_920_45156# 0.0109f
C4555 XA7.XA1.XA5.MN2.G a_14888_40228# 5.59e-19
C4556 XA2.XA4.MN0.D a_4808_42340# 9.25e-20
C4557 XA8.XA9.MN1.G a_21080_51140# 0.0222f
C4558 XA1.XA12.MP0.G VREF 0.0123f
C4559 AVDD a_8480_48676# 0.00129f
C4560 CK_SAMPLE a_18560_49380# 0.00139f
C4561 a_8480_51844# a_8480_51492# 0.0109f
C4562 a_18560_51844# XA7.XA8.MP0.D 0.0215f
C4563 XDAC1.XC0.XRES2.B XDAC1.XC64b<1>.XRES2.B 1.67e-19
C4564 li_9184_30036# li_9184_29616# 0.00411f
C4565 XA0.XA6.MP2.G li_9184_22656# 3.5e-20
C4566 XA20.XA2a.MN0.D a_12368_42340# 0.00768f
C4567 SARN XDAC2.XC1.XRES2.B 6.99f
C4568 XA0.XA1.XA5.MP1.D a_n232_43748# 2.16e-19
C4569 XA0.XA1.XA5.MN1.D a_920_43748# 2.16e-19
C4570 EN a_2288_43748# 0.166f
C4571 a_13520_44100# a_13520_43748# 0.0109f
C4572 XA20.XA3a.MN0.D XA1.XA1.XA1.MP1.D 0.0093f
C4573 AVDD a_23600_45508# 0.00149f
C4574 D<1> XA4.XA6.MP0.G 0.0317f
C4575 D<4> XA7.XA6.MP0.G 1.7e-19
C4576 SARN a_23600_48676# 0.156f
C4577 a_12368_51492# VREF 0.00396f
C4578 a_16040_50788# a_16040_50436# 0.0109f
C4579 D<3> XA6.XA6.MP0.G 0.121f
C4580 a_3440_50788# XA1.XA6.MP0.G 1.75e-20
C4581 D<2> XA5.XA6.MP0.G 0.026f
C4582 XDAC1.XC32a<0>.XRES8.B XDAC1.XC32a<0>.XRES2.B 0.44f
C4583 XDAC2.XC32a<0>.XRES8.B li_14804_14472# 9.91e-20
C4584 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES16.B 0.0483f
C4585 XA6.XA1.XA2.MP0.D a_16040_42340# 2.54e-19
C4586 XA5.XA1.XA4.MP1.D XA5.XA1.XA4.MN1.D 0.00918f
C4587 XA2.XA1.XA2.MP0.D a_5960_41988# 0.0219f
C4588 XA1.XA4.MN0.D li_9184_12216# 0.00504f
C4589 XA0.XA4.MN0.D XDAC1.XC64a<0>.XRES4.B 2.23e-21
C4590 EN XA5.XA1.XA1.MN0.S 0.139f
C4591 XA6.XA1.XA5.MN2.G a_11000_46564# 7.1e-20
C4592 XA5.XA1.XA5.MN2.G a_12368_46564# 7.1e-20
C4593 AVDD XA7.XA1.XA4.MP1.D 0.0913f
C4594 VREF a_5960_49028# 0.0647f
C4595 XA8.XA4.MN0.D a_21080_49380# 0.154f
C4596 a_22448_55364# XA20.XA12.MP0.G 0.00164f
C4597 a_22448_55012# a_23600_55012# 0.00133f
C4598 a_23600_55364# XA20.XA12.MP0.D 2.54e-19
C4599 AVDD a_22448_54660# 0.383f
C4600 SARP XDAC1.XC64b<1>.XRES16.B 55.3f
C4601 AVDD a_16040_40228# 0.467f
C4602 XA6.XA4.MN0.G a_14888_47268# 0.157f
C4603 D<7> a_3440_43748# 6.49e-19
C4604 XA4.XA1.XA5.MN2.G XA4.XA1.XA2.MP0.D 0.126f
C4605 XA20.XA3.MN0.D a_23600_45508# 0.0269f
C4606 VREF a_21080_45860# 0.0174f
C4607 XA2.XA11.MN1.G a_2288_52548# 7.25e-20
C4608 XA2.XA11.MP0.D XA2.XA10.MP0.D 0.00986f
C4609 a_8480_53252# a_9848_53252# 8.89e-19
C4610 AVDD a_22448_52196# 0.569f
C4611 a_11000_40228# a_12368_40228# 8.89e-19
C4612 XA8.XA7.MP0.G a_21080_41284# 0.0171f
C4613 XA5.XA3.MN0.G XA5.XA1.XA5.MN2.D 0.702f
C4614 D<8> a_920_45156# 0.0546f
C4615 XA2.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.D 0.0288f
C4616 XA5.XA6.MP0.G XA5.XA1.XA4.MN0.D 6.07e-19
C4617 a_12368_46212# a_12368_45860# 0.0109f
C4618 a_17408_52196# a_18560_52196# 0.00133f
C4619 a_17408_52900# XA8.XA1.XA5.MN2.G 1.06e-19
C4620 AVDD a_7328_49732# 0.359f
C4621 a_n232_52196# a_n232_51844# 0.0109f
C4622 a_7328_52196# XA3.XA7.MP0.D 0.0674f
C4623 CK_SAMPLE XA8.XA6.MN0.D 0.0433f
C4624 a_8408_334# a_9560_334# 0.00133f
C4625 a_13808_686# a_13808_334# 0.0109f
C4626 CK_SAMPLE_BSSW a_11000_334# 5.73e-19
C4627 XA7.XA1.XA5.MN2.D a_18560_43748# 0.00224f
C4628 XA20.XA2a.MN0.D a_19928_43044# 0.00118f
C4629 XA6.XA4.MN0.G a_14888_41636# 6.69e-20
C4630 a_5960_44452# a_5960_44100# 0.0109f
C4631 a_13520_44804# EN 7.78e-19
C4632 a_5960_51492# XA2.XA6.MP0.G 4.06e-20
C4633 XA20.XA9.MP0.D a_21080_48676# 5.7e-20
C4634 XA5.XA9.MN1.G XA5.XA4.MN0.D 0.00938f
C4635 AVDD a_11000_46564# 0.356f
C4636 a_13520_51140# a_13520_50788# 0.0109f
C4637 XA6.XA7.MP0.D a_14888_50084# 7.44e-20
C4638 XB2.XA3.MN1.D m3_16544_2420# 0.0137f
C4639 a_5960_43396# a_5960_43044# 0.0109f
C4640 XA20.XA2a.MN0.D a_18560_40580# 0.00123f
C4641 XA1.XA3.MN0.G a_3440_39876# 0.00646f
C4642 XA1.XA6.MP0.G XDAC2.XC64a<0>.XRES1B.B 0.00405f
C4643 AVDD XA3.XA1.XA5.MP0.D 0.159f
C4644 XA20.XA10.MN1.D a_23600_44452# 0.00405f
C4645 XA5.XA6.MP0.G a_13520_49380# 0.0547f
C4646 a_5960_50084# VREF 0.00382f
C4647 a_16040_50084# a_16040_49732# 0.0109f
C4648 a_2288_49732# a_3440_49732# 0.00133f
C4649 XA1.XA6.MP0.G a_3440_49028# 0.0137f
C4650 XA20.XA3a.MN0.G XA8.XA4.MN0.D 0.00217f
C4651 a_17408_42340# a_17408_41988# 0.0109f
C4652 D<8> XDAC2.XC128a<1>.XRES2.B 0.00406f
C4653 a_22448_48324# a_23600_48324# 0.00133f
C4654 D<1> a_18560_45156# 7.77e-19
C4655 AVDD XA0.XA1.XA1.MN0.D 0.0357f
C4656 XA5.XA4.MN0.D a_13520_46916# 0.00396f
C4657 D<5> a_7328_44804# 2.37e-19
C4658 XA8.XA1.XA5.MN2.G a_19928_44452# 5.11e-19
C4659 XA0.XA7.MP0.G a_3440_44100# 0.0693f
C4660 XA2.XA1.XA5.MN2.G a_2288_44100# 0.00556f
C4661 a_4808_48324# a_4808_47972# 0.0109f
C4662 XA6.XA11.MN1.G a_16040_53604# 0.0658f
C4663 AVDD a_19928_52900# 0.00166f
C4664 a_4808_40932# a_4808_40580# 0.0109f
C4665 XA6.XA1.XA1.MP1.D a_16040_40580# 0.00176f
C4666 XA1.XA1.XA1.MN0.D a_3440_40228# 0.00155f
C4667 XA6.XA1.XA1.MN0.S a_14888_39876# 2.54e-19
C4668 XA20.XA3a.MN0.D XA0.XA1.XA5.MN2.D 3.88e-19
C4669 XA0.XA11.MN1.G SAR_IP 0.374f
C4670 a_5960_46564# a_7328_46564# 8.89e-19
C4671 D<8> XA20.XA2a.MN0.D 0.244f
C4672 XA5.XA1.XA5.MN2.G a_9848_41988# 0.0684f
C4673 XA2.XA10.MP0.G a_5960_52196# 0.0441f
C4674 AVDD a_7328_50436# 0.416f
C4675 DONE a_19928_50788# 1.18e-19
C4676 a_9848_52548# XA4.XA9.MN1.G 0.0727f
C4677 CK_SAMPLE D<1> 0.0524f
C4678 XB2.XA4.MP0.D a_14960_2094# 0.0682f
C4679 SAR_IP a_11000_1390# 0.0597f
C4680 XB2.XA1.MP0.D XB2.XA3.MN1.D 4.9e-19
C4681 XB1.M1.G a_11000_1742# 0.00169f
C4682 XB2.M1.G XB2.XA0.MP0.D 0.303f
C4683 a_n232_44804# a_920_44804# 0.00133f
C4684 XA20.XA2a.MN0.D a_14888_43748# 4.48e-20
C4685 SARN li_14804_27780# 0.00103f
C4686 XA2.XA4.MN0.G XA2.XA1.XA4.MN0.D 0.00331f
C4687 XA20.XA3a.MN0.D XA7.XA1.XA4.MN1.D 0.0124f
C4688 XA3.XA1.XA5.MN2.D a_8480_44452# 0.153f
C4689 a_13520_45156# a_13520_44804# 0.0109f
C4690 XA3.XA1.XA5.MN2.G a_5960_51140# 0.077f
C4691 XA4.XA10.MP0.D VREF 0.0118f
C4692 XA3.XA9.MN1.G XA3.XA6.MP0.D 0.0618f
C4693 a_17408_51844# D<1> 1.25e-19
C4694 AVDD a_8480_47620# 0.00125f
C4695 SARN a_22448_50436# 6.57e-19
C4696 XB1.XA4.MP0.D XDAC1.XC1.XRES4.B 0.00738f
C4697 XDAC2.X16ab.XRES8.B XDAC2.X16ab.XRES2.B 0.44f
C4698 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES16.B 0.0483f
C4699 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES1A.B 0.00438f
C4700 XA20.XA2a.MN0.D a_2288_41284# 0.0685f
C4701 XA2.XA1.XA2.MP0.D XA2.XA1.XA5.MN0.D 0.056f
C4702 XA6.XA1.XA5.MN1.D a_14888_43396# 0.00176f
C4703 a_16040_43748# XA6.XA1.XA5.MP0.D 0.00176f
C4704 a_3440_43748# a_3440_43396# 0.0109f
C4705 D<6> li_9184_13248# 0.00504f
C4706 EN a_5960_43044# 0.141f
C4707 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES4.B 0.00405f
C4708 XA5.XA6.MP0.G XA7.XA6.MP0.G 0.318f
C4709 a_16040_50436# a_16040_50084# 0.0109f
C4710 XA20.XA10.MN1.D a_23600_45508# 0.00411f
C4711 XA20.XA9.MP0.D a_23600_46564# 0.00558f
C4712 XA1.XA6.MP0.G a_3440_50084# 6.4e-20
C4713 XA1.XA6.MP0.D a_2288_50084# 0.049f
C4714 AVDD a_22448_44452# 0.416f
C4715 SARN a_23600_47620# 0.0017f
C4716 XDAC2.XC64a<0>.XRES8.B XDAC2.XC1.XRES8.B 6.7e-19
C4717 li_14804_9768# li_14804_9156# 0.00271f
C4718 a_9848_42692# a_9848_42340# 0.0109f
C4719 XA8.XA1.XA4.MP1.D a_21080_42340# 0.00176f
C4720 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES2.B 0.00405f
C4721 XA8.XA4.MN0.D XA7.XA4.MN0.G 3.16e-20
C4722 XA7.XA4.MN0.D XA8.XA4.MN0.G 3.16e-20
C4723 AVDD a_8480_41988# 0.00125f
C4724 a_16040_49028# a_16040_48676# 0.0109f
C4725 VREF a_7328_47972# 0.0175f
C4726 XA2.XA4.MN0.D a_4808_47972# 0.0788f
C4727 XA8.XA1.XA5.MN2.G a_19928_45508# 9.01e-20
C4728 XA2.XA1.XA5.MN2.G XA2.XA1.XA5.MN2.D 0.0398f
C4729 a_5960_53956# a_7328_53956# 8.89e-19
C4730 a_19928_54308# a_19928_53956# 0.0109f
C4731 AVDD a_5960_53604# 0.383f
C4732 DONE XA8.XA11.MN1.G 0.00199f
C4733 a_7328_54308# XA4.XA11.MN1.G 8.3e-19
C4734 XA3.XA1.XA1.MP2.D a_7328_40932# 0.00176f
C4735 a_19928_41284# a_21080_41284# 0.00133f
C4736 SARP li_9184_17340# 0.00103f
C4737 XA6.XA4.MN0.G a_14888_46212# 0.0149f
C4738 XA7.XA1.XA5.MN2.G XA6.XA1.XA4.MN1.D 7.2e-19
C4739 XA6.XA1.XA5.MN2.G XA6.XA1.XA4.MP1.D 7.44e-19
C4740 a_11000_47268# a_11000_46916# 0.0109f
C4741 XA0.XA7.MP0.G a_n232_42692# 1.95e-19
C4742 VREF a_21080_44804# 0.069f
C4743 AVDD a_14960_2094# 0.362f
C4744 SARN a_23600_41988# 5.16e-19
C4745 AVDD a_2288_51140# 0.383f
C4746 XA20.XA10.MN1.D a_22448_52196# 1.97e-19
C4747 a_3440_53252# XA1.XA9.MN1.G 5.25e-19
C4748 a_14888_52900# a_16040_52900# 0.00133f
C4749 CK_SAMPLE XA7.XA8.MP0.D 3.93e-19
C4750 XA6.XA11.MN1.G XA5.XA7.MP0.D 4.87e-19
C4751 a_9560_3502# a_9560_3150# 0.0109f
C4752 XB1.XA2.MN0.G a_8408_3150# 0.0715f
C4753 XA20.XA3a.MN0.D XA3.XA1.XA5.MN0.D 0.0107f
C4754 a_8480_45508# XA3.XA1.XA5.MN2.D 0.0658f
C4755 XA4.XA4.MN0.G a_11000_43396# 8.07e-19
C4756 XA6.XA1.XA5.MN2.G a_14888_40228# 0.0709f
C4757 SARN XB2.XA3.MN1.D 8.04e-19
C4758 XA3.XA3.MN0.G a_7328_44100# 0.00245f
C4759 XA8.XA9.MN1.G a_19928_51140# 0.0469f
C4760 XA2.XA9.MN1.G XA2.XA6.MP2.D 0.0618f
C4761 XA2.XA11.MN1.G VREF 0.0162f
C4762 AVDD a_7328_48676# 0.356f
C4763 CK_SAMPLE a_17408_49380# 7.89e-19
C4764 a_17408_51844# XA7.XA8.MP0.D 0.0215f
C4765 XA1.XA7.MP0.D XA2.XA1.XA5.MN2.G 0.14f
C4766 XA7.XA7.MP0.D a_18560_51492# 0.126f
C4767 XA0.XA1.XA5.MN1.D a_n232_43748# 0.0494f
C4768 EN a_920_43748# 0.166f
C4769 D<5> XDAC1.X16ab.XRES16.B 0.00543f
C4770 XA20.XA3a.MN0.D XA0.XA1.XA1.MP1.D 0.0093f
C4771 XA8.XA1.XA5.MN2.D a_21080_43044# 1.88e-19
C4772 XA20.XA2a.MN0.D a_11000_42340# 0.00732f
C4773 AVDD a_22448_45508# 0.368f
C4774 a_11000_51492# VREF 0.00396f
C4775 D<3> XA5.XA6.MN0.D 0.00148f
C4776 a_2288_50436# a_3440_50436# 0.00133f
C4777 a_2288_50788# XA1.XA6.MP0.G 1.34e-19
C4778 XA2.XA1.XA2.MP0.D a_4808_41988# 0.0568f
C4779 XA6.XA1.XA2.MP0.D a_14888_42340# 0.095f
C4780 XA0.XA1.XA4.MP1.D a_920_42692# 0.049f
C4781 a_13520_43044# a_13520_42692# 0.0109f
C4782 XA5.XA1.XA5.MN2.G a_11000_46564# 0.00363f
C4783 a_8480_49380# a_9848_49380# 8.89e-19
C4784 AVDD XA6.XA1.XA4.MP1.D 0.0913f
C4785 XA4.XA6.MP0.G XA4.XA4.MN0.G 0.0415f
C4786 XA7.XA6.MP0.G a_18560_48324# 0.00295f
C4787 XA1.XA4.MN0.D a_3440_49028# 0.156f
C4788 XA8.XA4.MN0.D a_19928_49380# 0.155f
C4789 VREF a_4808_49028# 7.81e-19
C4790 a_23600_55364# a_23600_55012# 0.0109f
C4791 a_22448_55364# XA20.XA12.MP0.D 2.54e-19
C4792 AVDD XA20.XA12.MP0.G 1.64f
C4793 a_n232_41636# a_n232_41284# 0.0109f
C4794 a_11000_41636# XA4.XA1.XA1.MP2.D 0.00176f
C4795 AVDD a_14888_40228# 0.00131f
C4796 a_17408_47972# a_17408_47620# 0.0109f
C4797 a_3440_47620# a_4808_47620# 8.89e-19
C4798 D<7> a_2288_43748# 7.77e-20
C4799 XA3.XA1.XA5.MN2.G XA4.XA1.XA2.MP0.D 1.74e-19
C4800 XA4.XA1.XA5.MN2.G XA3.XA1.XA5.MN0.D 7.2e-19
C4801 XA5.XA4.MN0.D a_13520_45860# 5.88e-20
C4802 VREF a_19928_45860# 1.19e-19
C4803 a_19928_53604# XA8.XA10.MP0.D 1.17e-19
C4804 XA5.XA11.MN1.G XA5.XA10.MP0.G 0.0119f
C4805 CK_SAMPLE XA2.XA9.MN1.G 0.134f
C4806 XA8.XA12.MP0.G a_21080_52900# 1.28e-19
C4807 XA0.XA12.MP0.D a_3440_52548# 0.00103f
C4808 AVDD a_21080_52196# 0.37f
C4809 a_23600_40580# a_23600_40228# 0.0109f
C4810 XA1.XA6.MP0.G a_3440_42340# 7.76e-20
C4811 XA8.XA7.MP0.G a_19928_41284# 0.00527f
C4812 D<8> a_n232_45156# 0.083f
C4813 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MN0.D 0.0825f
C4814 XA8.XA4.MN0.G EN 0.0569f
C4815 XA2.XA4.MN0.G XA2.XA1.XA5.MP1.D 0.00138f
C4816 XA5.XA6.MP0.G XA5.XA1.XA4.MP0.D 9.97e-19
C4817 XA0.XA10.MP0.G XA0.XA7.MP0.G 2.18e-19
C4818 AVDD a_5960_49732# 0.359f
C4819 CK_SAMPLE XA8.XA6.MP0.G 0.00921f
C4820 CK_SAMPLE_BSSW a_9560_334# 0.0832f
C4821 SARN XDAC2.XC128a<1>.XRES2.B 6.99f
C4822 XA20.XA3a.MN0.D a_9848_41988# 0.00547f
C4823 a_17408_44452# a_18560_44452# 0.00133f
C4824 XA7.XA1.XA5.MN2.D a_17408_43748# 0.00388f
C4825 XA20.XA2a.MN0.D a_18560_43044# 1.43e-19
C4826 XA2.XA3.MN0.G a_4808_42692# 0.00335f
C4827 a_12368_44804# EN 3.4e-19
C4828 XA0.XA6.MP2.G li_9184_33096# 0.00508f
C4829 XA3.XA4.MN0.D a_8480_40580# 9.24e-20
C4830 AVDD a_9848_46564# 0.00125f
C4831 XA0.XA6.MP2.G a_920_50788# 0.161f
C4832 XA0.XA6.MN2.D a_n232_50788# 0.0488f
C4833 XA1.XA9.MN1.G a_3440_49380# 4.23e-20
C4834 XA7.XA9.MN1.G VREF 0.0732f
C4835 XDAC1.XC128b<2>.XRES1A.B XDAC1.XC128a<1>.XRES1B.B 0.617f
C4836 XB2.XA3.MN1.D m3_16472_2420# 0.0137f
C4837 a_17408_43396# a_18560_43396# 0.00133f
C4838 XA7.XA1.XA5.MP0.D a_17408_43044# 0.00176f
C4839 XA7.XA1.XA2.MP0.D a_18560_43044# 0.0292f
C4840 XA3.XA1.XA2.MP0.D XA3.XA1.XA4.MN1.D 0.056f
C4841 SARP a_23600_41988# 0.165f
C4842 EN XA8.XA1.XA4.MP0.D 0.0386f
C4843 XA0.XA4.MN0.D XDAC1.XC128b<2>.XRES4.B 0.00405f
C4844 XA0.XA6.MP0.G li_14804_12216# 1.85e-20
C4845 XA6.XA6.MP0.G XDAC2.XC32a<0>.XRES8.B 4.63e-20
C4846 AVDD XA3.XA1.XA2.MP0.D 0.263f
C4847 D<5> XA3.XA4.MN0.G 0.259f
C4848 SARN XA20.XA2a.MN0.D 0.00451f
C4849 XA20.XA10.MN1.D a_22448_44452# 1.87e-19
C4850 XA5.XA6.MP0.G a_12368_49380# 0.0781f
C4851 a_3440_50084# XA1.XA4.MN0.D 3.12e-20
C4852 XA1.XA6.MP0.G a_2288_49028# 0.0307f
C4853 a_3440_41988# a_4808_41988# 8.89e-19
C4854 D<1> a_17408_45156# 6.68e-19
C4855 a_13520_48324# XA5.XA4.MN0.G 0.0661f
C4856 AVDD a_23600_41284# 0.00183f
C4857 XA5.XA4.MN0.D a_12368_46916# 0.00245f
C4858 XA8.XA1.XA5.MN2.G a_18560_44452# 1.86e-19
C4859 XA0.XA7.MP0.G a_2288_44100# 7.1e-20
C4860 XA2.XA1.XA5.MN2.G a_920_44100# 7.1e-20
C4861 XA2.XA11.MN1.G XA0.XA11.MN1.G 1.54e-19
C4862 XA6.XA11.MN1.G a_14888_53604# 0.0709f
C4863 XA5.XA12.MP0.G a_13520_53604# 0.102f
C4864 AVDD a_18560_52900# 0.00166f
C4865 XA0.XA12.MP0.D XA1.XA11.MP0.D 0.0383f
C4866 XA0.XA12.MP0.G XA0.XA11.MP0.D 0.0612f
C4867 a_920_53604# a_2288_53604# 8.89e-19
C4868 a_16040_40932# a_17408_40932# 8.89e-19
C4869 XA6.XA1.XA1.MN0.D a_16040_40580# 8.3e-19
C4870 SARP XDAC1.XC1.XRES2.B 6.99f
C4871 XA20.XA3a.MN0.D a_23600_45508# 5.28e-19
C4872 XA0.XA11.MN1.G XB1.XA1.MN0.D 0.00904f
C4873 XA6.XA4.MN0.G a_16040_45156# 5.54e-19
C4874 XA6.XA3.MN0.G a_16040_46564# 0.155f
C4875 a_23600_46916# XA20.XA2a.MN0.D 7.42e-20
C4876 XA4.XA1.XA5.MN2.G a_9848_41988# 0.00407f
C4877 D<4> XA4.XA1.XA4.MP0.D 6.08e-19
C4878 XA2.XA4.MN0.D a_5960_43748# 9.14e-20
C4879 XA2.XA10.MP0.G a_4808_52196# 0.0131f
C4880 XA8.XA10.MP0.G XA8.XA9.MN0.D 0.106f
C4881 CK_SAMPLE XA6.XA6.MP2.D 3.06e-19
C4882 AVDD a_5960_50436# 0.416f
C4883 a_21080_52548# a_22448_52548# 8.89e-19
C4884 SAR_IP a_9560_1390# 0.00815f
C4885 XB1.XA4.MP0.D a_8408_1742# 0.015f
C4886 SAR_IN XB2.XA3.MN1.D 0.234f
C4887 XB2.XA1.MP0.D XB2.XA3.MN0.S 6.58e-19
C4888 a_9560_2094# a_11000_2094# 8e-19
C4889 XB1.M1.G a_9560_1742# 0.00285f
C4890 a_8408_2446# XB1.XA3.MN1.D 4.69e-19
C4891 a_9560_2446# XB1.XA3.MN0.S 1.03e-19
C4892 XA8.XA4.MN0.G a_21080_42692# 0.00224f
C4893 XA6.XA6.MP0.G a_16040_40932# 4.24e-19
C4894 XA5.XA3.MN0.G XA5.XA1.XA2.MP0.D 0.00212f
C4895 XA2.XA6.MP0.G a_5960_40580# 5.5e-19
C4896 XA20.XA3a.MN0.D XA7.XA1.XA4.MP1.D 0.0124f
C4897 XA3.XA1.XA5.MN2.D a_7328_44452# 0.158f
C4898 XA20.XA2a.MN0.D a_13520_43748# 2.91e-20
C4899 XA3.XA1.XA5.MN2.G a_4808_51140# 0.0661f
C4900 XA8.XA1.XA5.MN2.G XA8.XA7.MP0.G 0.0185f
C4901 XA3.XA10.MP0.D VREF 0.0118f
C4902 XA3.XA9.MN1.G XA3.XA6.MP0.G 0.0725f
C4903 XA5.XA7.MP0.D a_13520_50788# 3.29e-19
C4904 a_16040_51492# a_16040_51140# 0.0109f
C4905 AVDD a_7328_47620# 0.356f
C4906 XA20.XA2a.MN0.D a_920_41284# 0.0669f
C4907 XA3.XA3.MN0.G XA3.XA1.XA1.MN0.D 0.00142f
C4908 EN a_4808_43044# 6.46e-19
C4909 D<1> li_9184_15696# 0.00504f
C4910 D<3> XDAC1.XC32a<0>.XRES8.B 4.63e-20
C4911 XA20.XA10.MN1.D a_22448_45508# 1.78e-19
C4912 XA0.XA6.MP2.G a_920_49028# 0.00884f
C4913 D<4> a_11000_49380# 0.00891f
C4914 XA1.XA6.MP0.G a_2288_50084# 0.159f
C4915 AVDD a_21080_44452# 0.357f
C4916 D<8> XDAC2.XC64b<1>.XRES2.B 4.06e-21
C4917 XA8.XA1.XA2.MP0.D XA8.XA1.XA1.MN0.S 2.11e-19
C4918 a_21080_42692# XA8.XA1.XA4.MP0.D 0.00176f
C4919 XA7.XA6.MP0.G a_18560_47268# 1.38e-19
C4920 XA7.XA4.MN0.D XA7.XA4.MN0.G 0.707f
C4921 AVDD a_7328_41988# 0.386f
C4922 XA3.XA6.MP0.G a_8480_46916# 7.76e-20
C4923 a_2288_48676# a_3440_48676# 0.00133f
C4924 VREF a_5960_47972# 0.0175f
C4925 XA8.XA1.XA5.MN2.G a_18560_45508# 2.31e-19
C4926 XA2.XA1.XA5.MN2.G XA1.XA1.XA5.MN2.D 0.108f
C4927 AVDD a_4808_53604# 0.00166f
C4928 XA20.XA12.MP0.G XA20.XA10.MN1.D 2.01e-19
C4929 XA20.XA11.MN0.D XA8.XA11.MN1.G 0.00217f
C4930 XA20.XA12.MP0.D XA20.XA10.MN0.D 0.0093f
C4931 a_8480_54308# XA3.XA11.MN1.G 0.00123f
C4932 XA3.XA1.XA1.MN0.S a_7328_40932# 0.0271f
C4933 a_7328_41284# XA3.XA1.XA1.MP1.D 0.00176f
C4934 XA6.XA4.MN0.G a_13520_46212# 2.2e-19
C4935 XA5.XA4.MN0.G a_14888_46212# 2.2e-19
C4936 XA6.XA1.XA5.MN2.G XA6.XA1.XA4.MN1.D 0.0131f
C4937 a_22448_47268# a_23600_47268# 0.00133f
C4938 VREF a_19928_44804# 7.12e-19
C4939 AVDD a_13808_2094# 0.00154f
C4940 XA5.XA6.MP0.G XA5.XA1.XA5.MN1.D 7.41e-19
C4941 AVDD a_920_51140# 0.383f
C4942 XA1.XA10.MP0.D a_3440_52548# 0.00316f
C4943 a_3440_52900# XA1.XA10.MP0.G 0.0665f
C4944 XA7.XA10.MP0.D XA7.XA10.MP0.G 0.194f
C4945 CK_SAMPLE XA6.XA8.MP0.D 3.93e-19
C4946 XA2.XA11.MN1.G a_3440_51844# 1.13e-19
C4947 XA20.XA3a.MN0.D XA3.XA1.XA5.MP0.D 7.25e-19
C4948 a_17408_45508# a_18560_45508# 0.00133f
C4949 a_7328_45508# XA3.XA1.XA5.MN2.D 0.0675f
C4950 a_n232_45508# a_n232_45156# 0.0109f
C4951 XA20.XA2a.MN0.D SARP 0.0291f
C4952 XA4.XA4.MN0.G a_9848_43396# 0.0104f
C4953 XA6.XA1.XA5.MN2.G a_13520_40228# 1.34e-19
C4954 XA5.XA1.XA5.MN2.G a_14888_40228# 4.72e-19
C4955 SARN XB2.XA3.MN0.S 0.00201f
C4956 XA7.XA6.MP0.G a_18560_41636# 7.76e-20
C4957 XA1.XA4.MN0.D a_3440_42340# 9.24e-20
C4958 XA8.XA9.MN1.G a_18560_51140# 2.84e-19
C4959 AVDD a_5960_48676# 0.356f
C4960 CK_SAMPLE a_16040_49380# 7.89e-19
C4961 a_17408_52196# XA8.XA1.XA5.MN2.G 3.39e-19
C4962 a_7328_51844# a_7328_51492# 0.0109f
C4963 XA7.XA7.MP0.D a_17408_51492# 0.0877f
C4964 XA0.XA12.MP0.G VREF 0.0119f
C4965 XA2.XA9.MN1.G XA2.XA6.MN2.D 0.126f
C4966 XDAC2.XC0.XRES1A.B XDAC2.XC64b<1>.XRES1B.B 0.617f
C4967 XA0.XA6.MP2.G XDAC1.XC128b<2>.XRES1B.B 4.06e-21
C4968 a_12368_44100# a_12368_43748# 0.0109f
C4969 EN a_n232_43748# 0.0785f
C4970 a_n232_44100# XA0.XA1.XA2.MP0.D 2.92e-19
C4971 SARN li_14804_7512# 0.00103f
C4972 XA20.XA3a.MN0.D XA0.XA1.XA1.MN0.D 0.0616f
C4973 XA8.XA1.XA5.MN2.D a_19928_43044# 5.1e-20
C4974 XA20.XA2a.MN0.D a_9848_42340# 0.0843f
C4975 a_9848_44452# XA4.XA1.XA2.MP0.D 5.16e-20
C4976 XA4.XA1.XA5.MN1.D XA4.XA1.XA5.MP1.D 0.00918f
C4977 XA4.XA1.XA5.MN2.G a_7328_49732# 0.00457f
C4978 D<3> XA5.XA6.MP0.D 0.0323f
C4979 XA0.XA6.MP2.G a_920_50084# 0.0155f
C4980 a_14888_50788# a_14888_50436# 0.0109f
C4981 AVDD a_21080_45508# 0.359f
C4982 XDAC1.XC32a<0>.XRES8.B li_9184_14472# 9.91e-20
C4983 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES2.B 0.0307f
C4984 li_14804_15084# li_14804_14472# 0.00271f
C4985 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES16.B 0.0381f
C4986 XA0.XA1.XA4.MP1.D a_n232_42692# 2.16e-19
C4987 XA0.XA1.XA4.MN1.D a_920_42692# 2.16e-19
C4988 XA1.XA4.MN0.D XDAC1.XC64a<0>.XRES1B.B 0.00405f
C4989 XA0.XA4.MN0.D li_9184_12216# 1.85e-20
C4990 EN XA4.XA1.XA1.MN0.S 0.139f
C4991 AVDD XA6.XA1.XA4.MN1.D 0.00889f
C4992 XA7.XA6.MP0.G a_17408_48324# 0.00417f
C4993 XA1.XA4.MN0.D a_2288_49028# 0.154f
C4994 VREF a_3440_49028# 7.81e-19
C4995 XA1.XA6.MP0.G a_3440_47972# 6.28e-19
C4996 AVDD XA20.XA12.MP0.D 1.16f
C4997 SARP li_9184_27780# 0.00103f
C4998 a_22448_41636# a_23600_41636# 0.00133f
C4999 a_11000_41636# XA4.XA1.XA1.MN0.S 0.0694f
C5000 AVDD a_13520_40228# 0.00131f
C5001 XA5.XA4.MN0.G a_13520_47268# 0.157f
C5002 XA4.XA1.XA5.MN2.G XA3.XA1.XA5.MP0.D 0.00353f
C5003 XA20.XA10.MN1.D a_23600_41284# 0.00505f
C5004 VREF a_18560_45860# 1.19e-19
C5005 XA1.XA11.MP0.D XA1.XA10.MP0.D 0.00986f
C5006 XA5.XA11.MN1.G XA4.XA10.MP0.G 0.0024f
C5007 XA8.XA12.MP0.G a_19928_52900# 0.00258f
C5008 a_7328_53252# a_8480_53252# 0.00133f
C5009 XA0.XA12.MP0.D a_2288_52548# 0.00135f
C5010 AVDD a_19928_52196# 0.00154f
C5011 a_9848_40228# a_11000_40228# 0.00133f
C5012 XA20.XA3a.MN0.D a_22448_44452# 0.0064f
C5013 XA4.XA3.MN0.G XA4.XA1.XA5.MN2.D 0.702f
C5014 XA1.XA6.MP0.G a_2288_42340# 5.5e-19
C5015 XA8.XA1.XA5.MN2.G a_19928_41284# 0.0044f
C5016 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MP1.D 0.148f
C5017 XA0.XA7.MP0.G XA1.XA1.XA1.MN0.D 0.0326f
C5018 XA3.XA4.MN0.D a_8480_43044# 9.24e-20
C5019 XA2.XA4.MN0.G XA2.XA1.XA5.MN1.D 0.0242f
C5020 XA7.XA4.MN0.G EN 0.0578f
C5021 XA20.XA2a.MN0.D a_23600_45860# 0.0163f
C5022 a_11000_46212# a_11000_45860# 0.0109f
C5023 a_16040_52196# a_17408_52196# 8.89e-19
C5024 a_16040_52900# XA7.XA1.XA5.MN2.G 1.06e-19
C5025 AVDD a_4808_49732# 0.00159f
C5026 a_5960_52196# XA2.XA7.MP0.D 0.0658f
C5027 CK_SAMPLE XA7.XA6.MN0.D 0.0676f
C5028 XA4.XA9.MN0.D a_9848_51844# 0.00176f
C5029 XA4.XA9.MN1.G a_11000_51844# 6.57e-19
C5030 CK_SAMPLE_BSSW a_8408_334# 0.0663f
C5031 a_12368_686# a_12368_334# 0.0109f
C5032 XA20.XA3a.MN0.D a_8480_41988# 0.00547f
C5033 XA0.XA1.XA5.MN2.D XA0.XA1.XA2.MP0.D 4.72e-19
C5034 XA5.XA4.MN0.G a_13520_41636# 6.69e-20
C5035 XA1.XA3.MN0.G a_4808_42692# 4.4e-20
C5036 XA2.XA3.MN0.G a_3440_42692# 4.21e-19
C5037 a_4808_44452# a_4808_44100# 0.0109f
C5038 a_11000_44804# EN 3.4e-19
C5039 XA3.XA4.MN0.D a_7328_40580# 9.15e-20
C5040 D<5> D<2> 0.00204f
C5041 D<4> D<3> 5.83f
C5042 AVDD a_8480_46564# 0.00125f
C5043 a_12368_51140# a_12368_50788# 0.0109f
C5044 D<6> D<1> 0.0356f
C5045 XA1.XA9.MN1.G a_2288_49380# 2.54e-19
C5046 XA5.XA7.MP0.D a_13520_50084# 7.44e-20
C5047 XA4.XA1.XA5.MN2.G a_7328_50436# 0.0046f
C5048 XB2.XA3.MN1.D m3_26048_3300# 0.17f
C5049 EN XA8.XA1.XA4.MN0.D 3.17e-19
C5050 XA7.XA1.XA2.MP0.D a_17408_43044# 3.59e-19
C5051 XA3.XA1.XA2.MP0.D XA3.XA1.XA4.MP1.D 4.34e-19
C5052 a_4808_43396# a_4808_43044# 0.0109f
C5053 AVDD XA2.XA1.XA5.MP0.D 0.159f
C5054 D<2> a_16040_48324# 0.0164f
C5055 SARN a_23600_46564# 0.00206f
C5056 a_14888_50084# a_14888_49732# 0.0109f
C5057 a_920_49732# a_2288_49732# 8.89e-19
C5058 a_16040_42692# XA6.XA1.XA1.MN0.S 6.76e-20
C5059 a_16040_42340# a_16040_41988# 0.0109f
C5060 D<8> li_14804_17952# 0.00508f
C5061 XA3.XA6.MP0.G a_8480_45860# 7.76e-20
C5062 a_12368_48324# XA5.XA4.MN0.G 0.0674f
C5063 a_21080_48324# a_22448_48324# 8.89e-19
C5064 XA7.XA6.MP0.G a_18560_46212# 4.4e-19
C5065 AVDD a_22448_41284# 0.569f
C5066 VREF a_17408_46916# 0.0536f
C5067 XA8.XA1.XA5.MN2.G a_17408_44452# 0.00486f
C5068 XA7.XA1.XA5.MN2.G a_18560_44452# 5.11e-19
C5069 XA0.XA7.MP0.G a_920_44100# 0.00556f
C5070 a_3440_48324# a_3440_47972# 0.0109f
C5071 XA6.XA11.MN1.G a_13520_53604# 0.00787f
C5072 XA5.XA12.MP0.G a_12368_53604# 0.0877f
C5073 AVDD a_17408_52900# 0.387f
C5074 XA0.XA12.MP0.D XA0.XA11.MP0.D 0.00856f
C5075 XA0.XA12.MP0.G XA0.XA11.MN1.G 0.21f
C5076 XA6.XA1.XA1.MN0.D a_14888_40580# 0.035f
C5077 a_3440_40932# a_3440_40580# 0.0109f
C5078 XA20.XA3a.MN0.D a_22448_45508# 0.0049f
C5079 XA2.XA6.MP0.G a_5960_43044# 5.5e-19
C5080 XA0.XA11.MN1.G XB1.XA1.MP0.D 0.0452f
C5081 a_4808_46564# a_5960_46564# 0.00133f
C5082 XA6.XA6.MP0.G a_16040_43396# 5.5e-19
C5083 XA6.XA4.MN0.G a_14888_45156# 0.00865f
C5084 XA6.XA3.MN0.G a_14888_46564# 0.156f
C5085 a_23600_46916# a_23600_46564# 0.0109f
C5086 XA0.XA6.MP2.G a_920_42340# 7.76e-20
C5087 XA4.XA1.XA5.MN2.G a_8480_41988# 0.0673f
C5088 D<4> XA4.XA1.XA4.MN0.D 0.00144f
C5089 XA2.XA4.MN0.D a_4808_43748# 9.25e-20
C5090 VREF a_7328_43748# 8.43e-19
C5091 XA8.XA10.MP0.G XA8.XA9.MN1.G 0.202f
C5092 a_8480_52548# XA3.XA9.MN0.D 0.00176f
C5093 CK_SAMPLE XA6.XA6.MN2.D 0.0389f
C5094 AVDD a_4808_50436# 0.00154f
C5095 XB1.XA1.MN0.D a_9560_1390# 3.62e-20
C5096 XB2.XA1.MN0.D XB2.XA3.MN1.D 2.08e-19
C5097 XB1.XA4.MN0.D XB1.XA0.MP0.D 0.012f
C5098 XB1.M1.G a_8408_1742# 0.0315f
C5099 SAR_IP a_8408_1390# 0.00155f
C5100 SAR_IN XB2.XA3.MN0.S 0.0903f
C5101 XB2.XA4.MN0.D a_13808_2094# 0.0492f
C5102 XB2.M1.G a_14960_2094# 0.0998f
C5103 XA1.XA4.MN0.G XA1.XA1.XA4.MN0.D 0.00331f
C5104 XA8.XA4.MN0.G a_19928_42692# 0.0049f
C5105 XA6.XA6.MP0.G a_14888_40932# 3.97e-20
C5106 D<1> a_19928_39876# 1.26e-19
C5107 SARN XDAC2.XC64b<1>.XRES2.B 6.99f
C5108 XA2.XA6.MP0.G a_4808_40580# 7.76e-20
C5109 XA20.XA3a.MN0.D XA6.XA1.XA4.MP1.D 0.0124f
C5110 a_12368_45156# a_12368_44804# 0.0109f
C5111 XA2.XA10.MP0.D VREF 0.0118f
C5112 a_2288_51492# D<7> 2.41e-19
C5113 AVDD a_5960_47620# 0.356f
C5114 XDAC1.X16ab.XRES8.B XDAC1.X16ab.XRES2.B 0.44f
C5115 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES16.B 0.0483f
C5116 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES1A.B 0.00438f
C5117 XDAC2.X16ab.XRES8.B li_14804_24912# 9.91e-20
C5118 XA20.XA2a.MN0.D a_n232_41284# 0.0895f
C5119 XA5.XA1.XA5.MN1.D a_13520_43396# 0.00176f
C5120 a_14888_43748# XA6.XA1.XA5.MN0.D 0.00176f
C5121 a_2288_43748# a_2288_43396# 0.0109f
C5122 D<6> XDAC1.XC32a<0>.XRES16.B 0.0186f
C5123 D<4> li_9184_14472# 0.00504f
C5124 EN a_3440_43044# 5.26e-19
C5125 XA0.XA6.MP0.G li_14804_22656# 0.00504f
C5126 a_14888_50436# a_14888_50084# 0.0109f
C5127 XA0.XA6.MP2.G a_n232_49028# 5.7e-19
C5128 XA4.XA1.XA5.MN2.G a_7328_48676# 0.00363f
C5129 D<4> a_9848_49380# 5.91e-19
C5130 a_2288_50788# VREF 0.00345f
C5131 AVDD a_19928_44452# 0.00154f
C5132 li_9184_9768# li_9184_9156# 0.00271f
C5133 XDAC1.XC64a<0>.XRES8.B XDAC1.XC1.XRES8.B 6.7e-19
C5134 EN a_2288_40580# 0.0731f
C5135 XA1.XA3.MN0.G li_14804_28392# 0.00504f
C5136 XA4.XA1.XA2.MP0.D a_11000_41284# 1.07e-19
C5137 XA3.XA1.XA4.MP0.D XA3.XA1.XA4.MN0.D 0.00918f
C5138 XA8.XA1.XA4.MN1.D a_19928_42340# 0.00176f
C5139 a_8480_42692# a_8480_42340# 0.0109f
C5140 XA7.XA6.MP0.G a_17408_47268# 5.95e-19
C5141 XA3.XA6.MP0.G a_7328_46916# 5.5e-19
C5142 a_14888_49028# a_14888_48676# 0.0109f
C5143 XA1.XA4.MN0.D a_3440_47972# 0.0788f
C5144 VREF a_4808_47972# 7.39e-19
C5145 XA8.XA1.XA5.MN2.G a_17408_45508# 0.00595f
C5146 XA7.XA1.XA5.MN2.G a_18560_45508# 9.01e-20
C5147 XA0.XA7.MP0.G XA1.XA1.XA5.MN2.D 0.0405f
C5148 XA2.XA1.XA5.MN2.G XA0.XA1.XA5.MN2.D 6.95e-19
C5149 AVDD a_5960_41988# 0.386f
C5150 a_4808_53956# a_5960_53956# 0.00133f
C5151 a_18560_54308# a_18560_53956# 0.0109f
C5152 AVDD a_3440_53604# 0.00166f
C5153 XA20.XA12.MP0.D XA20.XA10.MN1.D 0.125f
C5154 XA20.XA12.MP0.G XA8.XA12.MP0.G 0.124f
C5155 a_7328_54308# XA3.XA11.MN1.G 8.45e-19
C5156 XA7.XA1.XA1.MP2.D XA7.XA1.XA1.MP1.D 0.0488f
C5157 XA7.XA1.XA1.MN0.S XA7.XA1.XA1.MN0.D 0.0743f
C5158 a_18560_41284# a_19928_41284# 8.89e-19
C5159 SARP XDAC1.XC128a<1>.XRES2.B 6.99f
C5160 XA5.XA4.MN0.G a_13520_46212# 0.0149f
C5161 XA20.XA3.MN6.D a_22448_44100# 0.0672f
C5162 XA20.XA3a.MN0.G a_23600_44100# 8.29e-20
C5163 XA6.XA1.XA5.MN2.G XA5.XA1.XA4.MN1.D 7.2e-19
C5164 a_9848_47268# a_9848_46916# 0.0109f
C5165 VREF a_18560_44804# 7.12e-19
C5166 XA5.XA6.MP0.G XA5.XA1.XA5.MP1.D 0.00121f
C5167 AVDD a_n232_51140# 0.00166f
C5168 XA1.XA10.MP0.D a_2288_52548# 0.00224f
C5169 a_13520_52900# a_14888_52900# 8.89e-19
C5170 a_2288_52900# XA1.XA10.MP0.G 0.0674f
C5171 CK_SAMPLE XA5.XA8.MP0.D 3.93e-19
C5172 XA5.XA11.MN1.G XA5.XA7.MP0.D 0.00283f
C5173 a_9560_3502# XB1.XA2.MN0.G 0.0658f
C5174 a_8408_3502# a_8408_3150# 0.0109f
C5175 XA20.XA3a.MN0.D XA3.XA1.XA2.MP0.D 0.199f
C5176 XA20.XA2a.MN0.D a_23600_44804# 0.00301f
C5177 D<3> a_13520_40932# 5.26e-19
C5178 XA3.XA6.MP0.G XA3.XA1.XA1.MN0.S 0.0123f
C5179 D<7> a_3440_40580# 5.26e-19
C5180 XA5.XA1.XA5.MN2.G a_13520_40228# 0.0825f
C5181 XA6.XA1.XA5.MN2.G a_12368_40228# 0.00255f
C5182 XA7.XA6.MP0.G a_17408_41636# 5.5e-19
C5183 XA1.XA4.MN0.D a_2288_42340# 9.15e-20
C5184 XA2.XA3.MN0.G a_5960_44100# 0.00245f
C5185 AVDD a_4808_48676# 0.00129f
C5186 CK_SAMPLE a_14888_49380# 0.00139f
C5187 XA7.XA9.MN1.G a_19928_51140# 2.84e-19
C5188 a_16040_51844# XA6.XA8.MP0.D 0.0215f
C5189 XA0.XA7.MP0.D XA0.XA7.MP0.G 0.14f
C5190 XA0.XA12.MP0.D VREF 0.39f
C5191 XA2.XA9.MN1.G D<6> 0.0378f
C5192 D<5> li_9184_24300# 0.00504f
C5193 EN XA8.XA1.XA5.MP1.D 0.0544f
C5194 XA20.XA2a.MN0.D a_8480_42340# 0.0848f
C5195 a_19928_44804# XA8.XA1.XA2.MP0.D 2.6e-20
C5196 XA3.XA1.XA5.MN2.G a_7328_49732# 7.1e-20
C5197 XA4.XA1.XA5.MN2.G a_5960_49732# 7.1e-20
C5198 D<3> XA5.XA6.MP0.G 2.11f
C5199 XA0.XA6.MP2.G a_n232_50084# 5.7e-19
C5200 D<5> XA7.XA6.MP0.G 4.27e-19
C5201 D<2> XA4.XA6.MP0.G 0.026f
C5202 a_920_50436# a_2288_50436# 8.89e-19
C5203 D<4> XA6.XA6.MP0.G 2.33e-19
C5204 D<1> XA3.XA6.MP0.G 0.0345f
C5205 AVDD a_19928_45508# 0.00166f
C5206 XA0.XA1.XA4.MN1.D a_n232_42692# 0.0474f
C5207 a_12368_43044# a_12368_42692# 0.0109f
C5208 a_7328_49380# a_8480_49380# 0.00133f
C5209 D<6> a_5960_46916# 0.0185f
C5210 AVDD XA5.XA1.XA4.MN1.D 0.00889f
C5211 VREF a_2288_49028# 0.0647f
C5212 XA7.XA4.MN0.D a_18560_49380# 0.155f
C5213 D<2> a_16040_47268# 0.0148f
C5214 XA1.XA6.MP0.G a_2288_47972# 8.92e-19
C5215 a_22448_55364# a_22448_55012# 0.0109f
C5216 AVDD a_23600_55012# 0.00166f
C5217 a_9848_41636# XA4.XA1.XA1.MN0.S 0.0674f
C5218 a_16040_47972# a_16040_47620# 0.0109f
C5219 XA3.XA6.MP0.G a_8480_44804# 7.76e-20
C5220 XA5.XA4.MN0.G a_12368_47268# 0.155f
C5221 a_2288_47620# a_3440_47620# 0.00133f
C5222 XA4.XA1.XA5.MN2.G XA3.XA1.XA2.MP0.D 0.146f
C5223 D<4> XA4.XA1.XA5.MP1.D 7.42e-19
C5224 XA20.XA10.MN1.D a_22448_41284# 1.97e-19
C5225 VREF a_17408_45860# 0.0178f
C5226 AVDD a_12368_40228# 0.464f
C5227 a_18560_53604# XA7.XA10.MP0.D 1.17e-19
C5228 XA7.XA11.MP0.D a_17408_53252# 0.0494f
C5229 CK_SAMPLE XA1.XA9.MN1.G 0.135f
C5230 XA0.XA12.MP0.D a_920_52548# 9.29e-19
C5231 AVDD a_18560_52196# 0.00154f
C5232 a_22448_40580# a_22448_40228# 0.0109f
C5233 XA20.XA3a.MN0.D a_21080_44452# 3.15e-19
C5234 XA3.XA3.MN0.G XA4.XA1.XA5.MN2.D 0.00909f
C5235 XA8.XA1.XA5.MN2.G a_18560_41284# 0.00733f
C5236 XA0.XA7.MP0.G XA1.XA1.XA1.MP1.D 6.68e-19
C5237 XA3.XA4.MN0.D a_7328_43044# 9.15e-20
C5238 XA6.XA4.MN0.G EN 0.0579f
C5239 D<2> a_16040_41636# 7.76e-20
C5240 XA20.XA2a.MN0.D a_22448_45860# 0.00531f
C5241 a_22448_46212# a_23600_46212# 0.00133f
C5242 XA6.XA10.MP0.G a_14888_51492# 6.8e-20
C5243 AVDD a_3440_49732# 0.00159f
C5244 CK_SAMPLE XA7.XA6.MP0.D 0.0278f
C5245 XA8.XA9.MN0.D XA8.XA7.MP0.D 0.00986f
C5246 a_4808_52196# XA2.XA7.MP0.D 0.0678f
C5247 XA4.XA9.MN1.G a_9848_51844# 0.0164f
C5248 SARN li_14804_17952# 0.00103f
C5249 a_16040_44452# a_17408_44452# 8.89e-19
C5250 XA6.XA1.XA5.MN2.D a_16040_43748# 0.00388f
C5251 XA1.XA3.MN0.G a_3440_42692# 0.00343f
C5252 a_9848_44804# EN 7.78e-19
C5253 XA0.XA6.MP2.G XDAC1.XC0.XRES1B.B 0.00406f
C5254 XA8.XA9.MN1.G a_21080_49732# 0.0215f
C5255 XA4.XA9.MN1.G XA4.XA4.MN0.D 0.00938f
C5256 AVDD a_7328_46564# 0.356f
C5257 D<4> XA4.XA6.MP2.D 0.0399f
C5258 XA6.XA9.MN1.G VREF 0.0732f
C5259 XA4.XA1.XA5.MN2.G a_5960_50436# 7.1e-20
C5260 XA3.XA1.XA5.MN2.G a_7328_50436# 7.1e-20
C5261 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128a<1>.XRES8.B 6.7e-19
C5262 XB2.XA3.MN1.D m3_25976_3300# 0.0634f
C5263 li_14804_20208# li_14804_19596# 0.00271f
C5264 EN XA7.XA1.XA4.MN0.D 3.17e-19
C5265 XA0.XA4.MN0.D li_9184_22656# 0.00504f
C5266 XA0.XA6.MP0.G XDAC2.XC64a<0>.XRES1B.B 2.23e-21
C5267 XA1.XA6.MP0.G XDAC2.XC32a<0>.XRES1A.A 0.0216f
C5268 XA20.XA2a.MN0.D a_14888_40580# 0.00138f
C5269 a_16040_43396# a_17408_43396# 8.89e-19
C5270 D<2> a_14888_48324# 6.53e-19
C5271 a_2288_50084# VREF 0.00382f
C5272 XA0.XA6.MP2.G a_920_47972# 0.0147f
C5273 XA8.XA6.MP0.G XA8.XA4.MN0.D 0.631f
C5274 XA4.XA1.XA5.MN2.G a_7328_47620# 0.00363f
C5275 AVDD XA2.XA1.XA5.MN0.D 0.00889f
C5276 SARP XB1.XA3.MN1.D 8.04e-19
C5277 a_2288_41988# a_3440_41988# 0.00133f
C5278 XA3.XA6.MP0.G a_7328_45860# 5.5e-19
C5279 XA7.XA6.MP0.G a_17408_46212# 5.5e-19
C5280 AVDD a_21080_41284# 0.361f
C5281 VREF a_16040_46916# 0.0536f
C5282 XA4.XA4.MN0.D a_11000_46916# 0.00245f
C5283 XA7.XA1.XA5.MN2.G a_17408_44452# 7.1e-20
C5284 XA8.XA1.XA5.MN2.G a_16040_44452# 7.1e-20
C5285 XA0.XA7.MP0.G a_n232_44100# 2.31e-19
C5286 XA6.XA11.MN1.G a_12368_53604# 0.00979f
C5287 AVDD a_16040_52900# 0.387f
C5288 XA0.XA12.MP0.D XA0.XA11.MN1.G 0.0251f
C5289 a_n232_53604# a_920_53604# 0.00133f
C5290 SARP li_9184_7512# 0.00103f
C5291 XA5.XA1.XA1.MN0.S a_13520_39876# 2.54e-19
C5292 a_14888_40932# a_16040_40932# 0.00133f
C5293 XA20.XA3a.MN0.D a_21080_45508# 7.22e-19
C5294 XA2.XA6.MP0.G a_4808_43044# 7.76e-20
C5295 XA6.XA6.MP0.G a_14888_43396# 7.76e-20
C5296 XA6.XA4.MN0.G a_13520_45156# 2.2e-19
C5297 XA5.XA4.MN0.G a_14888_45156# 2.2e-19
C5298 XA0.XA6.MP2.G a_n232_42340# 6.49e-19
C5299 XA3.XA1.XA5.MN2.G a_8480_41988# 0.0039f
C5300 XA4.XA1.XA5.MN2.G a_7328_41988# 0.0734f
C5301 VREF a_5960_43748# 8.43e-19
C5302 XA1.XA10.MP0.G a_3440_52196# 0.0131f
C5303 a_8480_52548# XA3.XA9.MN1.G 0.0711f
C5304 CK_SAMPLE D<2> 0.0523f
C5305 AVDD a_3440_50436# 0.00154f
C5306 a_19928_52548# a_21080_52548# 0.00133f
C5307 XB1.XA1.MP0.D a_9560_1390# 5.87e-20
C5308 a_8408_2094# a_9560_2094# 0.00133f
C5309 XB2.XA1.MN0.D XB2.XA3.MN0.S 0.00304f
C5310 XB1.XA4.MP0.D XB1.XA0.MP0.D 0.134f
C5311 XB2.M1.G a_13808_2094# 0.0193f
C5312 D<1> a_18560_39876# 0.00212f
C5313 XA20.XA3a.MN0.D XA6.XA1.XA4.MN1.D 0.0124f
C5314 XA2.XA1.XA5.MN2.D a_5960_44452# 0.158f
C5315 AVDD a_4808_47620# 0.00125f
C5316 XA7.XA1.XA5.MN2.G XA8.XA1.XA5.MN2.G 1.58f
C5317 XA1.XA10.MP0.D VREF 0.0118f
C5318 XA2.XA1.XA5.MN2.G a_3440_51140# 0.0677f
C5319 a_14888_51492# a_14888_51140# 0.0109f
C5320 XA8.XA9.MN1.G a_21080_50436# 7.76e-19
C5321 XA3.XA6.MP0.G XDAC2.X16ab.XRES16.B 0.00136f
C5322 XA20.XA2a.MN0.D XA8.XA1.XA1.MP2.D 0.0103f
C5323 a_14888_43748# XA6.XA1.XA2.MP0.D 0.0702f
C5324 D<3> li_9184_15084# 0.00504f
C5325 EN a_2288_43044# 0.141f
C5326 D<1> XDAC1.XC32a<0>.XRES1B.B 0.00405f
C5327 XA3.XA1.XA5.MN2.G a_7328_48676# 7.1e-20
C5328 XA4.XA1.XA5.MN2.G a_5960_48676# 7.1e-20
C5329 XA0.XA6.MP0.D a_920_50084# 0.049f
C5330 a_920_50788# VREF 0.00345f
C5331 D<1> XA7.XA4.MN0.D 0.203f
C5332 XA4.XA6.MP0.G XA7.XA6.MP0.G 0.0907f
C5333 XA5.XA6.MP0.G XA6.XA6.MP0.G 6.58f
C5334 AVDD a_18560_44452# 0.00125f
C5335 EN a_920_40580# 0.0717f
C5336 D<8> li_14804_28392# 3.5e-20
C5337 a_19928_42692# XA8.XA1.XA4.MN0.D 0.00176f
C5338 D<2> a_16040_46212# 0.0202f
C5339 XA6.XA4.MN0.D XA6.XA4.MN0.G 0.707f
C5340 a_920_48676# a_2288_48676# 8.89e-19
C5341 XA1.XA4.MN0.D a_2288_47972# 0.0546f
C5342 VREF a_3440_47972# 7.39e-19
C5343 D<6> a_5960_45860# 0.0774f
C5344 XA7.XA1.XA5.MN2.G a_17408_45508# 7.1e-20
C5345 XA8.XA1.XA5.MN2.G a_16040_45508# 7.1e-20
C5346 XA0.XA7.MP0.G XA0.XA1.XA5.MN2.D 0.108f
C5347 AVDD a_4808_41988# 0.00125f
C5348 AVDD a_2288_53604# 0.383f
C5349 a_23600_55012# XA20.XA10.MN1.D 1.44e-19
C5350 XA20.XA12.MP0.D XA8.XA12.MP0.G 0.00217f
C5351 a_5960_54308# XA3.XA11.MN1.G 0.00177f
C5352 XA7.XA1.XA1.MN0.S XA7.XA1.XA1.MP1.D 0.0615f
C5353 XA2.XA1.XA1.MP2.D a_5960_40932# 0.00176f
C5354 a_5960_41284# XA2.XA1.XA1.MP1.D 0.00176f
C5355 XA5.XA4.MN0.G a_12368_46212# 3.46e-19
C5356 XA20.XA3a.MN0.G a_22448_44100# 0.0632f
C5357 XA1.XA6.MP0.G a_3440_43748# 7.76e-20
C5358 XA6.XA1.XA5.MN2.G XA5.XA1.XA4.MP1.D 0.00353f
C5359 XA5.XA1.XA5.MN2.G XA5.XA1.XA4.MN1.D 0.0131f
C5360 D<7> a_3440_43044# 6.49e-19
C5361 a_21080_47268# a_22448_47268# 8.89e-19
C5362 VREF a_17408_44804# 0.0691f
C5363 D<3> a_13520_43396# 6.49e-19
C5364 AVDD XA8.XA7.MP0.G 5.21f
C5365 XA6.XA10.MP0.D XA6.XA10.MP0.G 0.194f
C5366 CK_SAMPLE XA4.XA8.MP0.D 3.93e-19
C5367 XA0.XA12.MP0.D a_3440_51844# 3.12e-19
C5368 XA5.XA11.MN1.G XA4.XA7.MP0.D 8.25e-19
C5369 a_19928_53604# XA8.XA9.MN1.G 7.36e-20
C5370 a_8408_3502# XB1.XA2.MN0.G 0.0955f
C5371 XA20.XA3a.MN0.D XA2.XA1.XA5.MP0.D 7.08e-19
C5372 a_16040_45508# a_17408_45508# 8.89e-19
C5373 a_5960_45508# XA2.XA1.XA5.MN2.D 0.0659f
C5374 XA20.XA2a.MN0.D a_22448_44804# 0.00157f
C5375 D<3> a_12368_40932# 4.18e-20
C5376 XA3.XA4.MN0.G a_8480_43396# 0.0104f
C5377 D<7> a_2288_40580# 4.18e-20
C5378 XA5.XA1.XA5.MN2.G a_12368_40228# 0.0128f
C5379 SARN XB1.XA3.MN0.S 9.84e-21
C5380 XA2.XA3.MN0.G a_4808_44100# 0.00768f
C5381 AVDD a_3440_48676# 0.00129f
C5382 CK_SAMPLE a_13520_49380# 0.00139f
C5383 XA7.XA9.MN1.G a_18560_51140# 0.0469f
C5384 a_16040_52196# XA7.XA1.XA5.MN2.G 3.39e-19
C5385 a_5960_51844# a_5960_51492# 0.0109f
C5386 a_14888_51844# XA6.XA8.MP0.D 0.0215f
C5387 XA6.XA7.MP0.D a_16040_51492# 0.0893f
C5388 XDAC1.XC0.XRES1A.B XDAC1.XC64b<1>.XRES1B.B 0.617f
C5389 SARN XDAC2.XC1.XRES8.B 27.7f
C5390 a_11000_44100# a_11000_43748# 0.0109f
C5391 EN XA8.XA1.XA5.MN1.D 0.0157f
C5392 XA7.XA1.XA5.MN2.D a_18560_43044# 5.1e-20
C5393 XA20.XA2a.MN0.D a_7328_42340# 0.00768f
C5394 D<6> XDAC1.X16ab.XRES16.B 9.19e-20
C5395 XA0.XA6.MP2.G li_9184_23076# 3.5e-20
C5396 a_7328_51492# VREF 0.00396f
C5397 XA3.XA1.XA5.MN2.G a_5960_49732# 0.00457f
C5398 XA8.XA7.MP0.G XA20.XA3.MN0.D 8.03e-19
C5399 a_13520_50788# a_13520_50436# 0.0109f
C5400 AVDD a_18560_45508# 0.00131f
C5401 li_9184_15084# li_9184_14472# 0.00271f
C5402 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES2.B 0.0307f
C5403 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES16.B 0.0381f
C5404 XA4.XA1.XA4.MN1.D XA4.XA1.XA4.MP1.D 0.00918f
C5405 XA0.XA4.MN0.D XDAC1.XC64a<0>.XRES1B.B 2.23e-21
C5406 EN XA3.XA1.XA1.MN0.S 0.139f
C5407 D<6> a_4808_46916# 0.00249f
C5408 AVDD XA5.XA1.XA4.MP1.D 0.0913f
C5409 VREF a_920_49028# 0.0647f
C5410 XA7.XA4.MN0.D a_17408_49380# 0.154f
C5411 D<2> a_14888_47268# 3.18e-19
C5412 a_22448_55364# a_23600_55364# 0.00133f
C5413 AVDD a_22448_55012# 0.467f
C5414 SARP XDAC1.XC64b<1>.XRES2.B 6.99f
C5415 a_21080_41636# a_22448_41636# 8.89e-19
C5416 D<1> EN 0.0683f
C5417 XA3.XA6.MP0.G a_7328_44804# 5.5e-19
C5418 XA3.XA1.XA5.MN2.G XA3.XA1.XA2.MP0.D 0.126f
C5419 D<4> XA4.XA1.XA5.MN1.D 0.00185f
C5420 XA7.XA6.MP0.G a_18560_45156# 7.76e-20
C5421 VREF a_16040_45860# 0.0178f
C5422 AVDD a_11000_40228# 0.467f
C5423 XA0.XA11.MP0.D XA0.XA10.MP0.D 0.00986f
C5424 XA7.XA12.MP0.G a_18560_52900# 0.00258f
C5425 XA8.XA11.MN1.G a_19928_52900# 7.39e-19
C5426 a_5960_53252# a_7328_53252# 8.89e-19
C5427 a_n232_53956# XA0.XA9.MN1.G 7.37e-20
C5428 AVDD a_17408_52196# 0.37f
C5429 XA4.XA11.MN1.G XA4.XA10.MP0.G 7.66e-19
C5430 a_8480_40228# a_9848_40228# 8.89e-19
C5431 XA3.XA3.MN0.G XA3.XA1.XA5.MN2.D 0.755f
C5432 XA8.XA1.XA5.MN2.G a_17408_41284# 0.0169f
C5433 XA7.XA1.XA5.MN2.G a_18560_41284# 0.00392f
C5434 D<6> XA2.XA1.XA1.MN0.S 0.0149f
C5435 XA0.XA7.MP0.G XA0.XA1.XA1.MP1.D 0.144f
C5436 XA1.XA4.MN0.G XA1.XA1.XA5.MN1.D 0.0242f
C5437 XA5.XA4.MN0.G EN 0.0578f
C5438 XA8.XA4.MN0.G a_21080_44100# 6.11e-19
C5439 D<2> a_14888_41636# 6.49e-19
C5440 a_9848_46212# a_9848_45860# 0.0109f
C5441 AVDD a_2288_49732# 0.359f
C5442 CK_SAMPLE XA7.XA6.MP0.G 0.0463f
C5443 XA8.XA9.MN1.G XA8.XA7.MP0.D 0.274f
C5444 a_14888_52196# a_16040_52196# 0.00133f
C5445 XA4.XA9.MN1.G a_8480_51844# 2.2e-19
C5446 a_14960_686# CK_SAMPLE_BSSW 0.0658f
C5447 a_11000_686# a_11000_334# 0.0109f
C5448 XA6.XA1.XA5.MN2.D a_14888_43748# 0.00224f
C5449 XA20.XA2a.MN0.D a_14888_43044# 1.43e-19
C5450 a_3440_44452# a_3440_44100# 0.0109f
C5451 a_8480_44804# EN 7.78e-19
C5452 XA2.XA4.MN0.D a_5960_40580# 9.14e-20
C5453 XA8.XA9.MN1.G a_19928_49732# 0.00119f
C5454 AVDD a_5960_46564# 0.356f
C5455 a_11000_51140# a_11000_50788# 0.0109f
C5456 D<4> XA4.XA6.MN2.D 1.59e-19
C5457 XA3.XA1.XA5.MN2.G a_5960_50436# 0.0046f
C5458 XB2.XA3.MN1.D m3_16544_3476# 0.0137f
C5459 D<8> a_n232_39876# 0.00627f
C5460 EN XA7.XA1.XA4.MP0.D 0.0386f
C5461 XA5.XA6.MP0.G XDAC2.XC32a<0>.XRES8.B 4.63e-20
C5462 XA7.XA6.MP0.G li_14804_15696# 0.00504f
C5463 XA20.XA2a.MN0.D a_13520_40580# 0.00123f
C5464 XA6.XA1.XA5.MP0.D a_16040_43044# 0.00176f
C5465 a_3440_43396# a_3440_43044# 0.0109f
C5466 a_n232_49732# a_920_49732# 0.00133f
C5467 a_13520_50084# a_13520_49732# 0.0109f
C5468 a_920_50084# VREF 0.00382f
C5469 XA0.XA6.MP2.G a_n232_47972# 5.43e-19
C5470 XA3.XA1.XA5.MN2.G a_7328_47620# 7.1e-20
C5471 XA4.XA1.XA5.MN2.G a_5960_47620# 7.1e-20
C5472 AVDD XA2.XA1.XA2.MP0.D 0.263f
C5473 SARP XB1.XA3.MN0.S 0.00202f
C5474 a_14888_42340# a_14888_41988# 0.0109f
C5475 D<8> XDAC2.XC128a<1>.XRES8.B 0.00688f
C5476 D<6> a_5960_44804# 2.36e-19
C5477 a_11000_48324# XA4.XA4.MN0.G 0.0658f
C5478 a_19928_48324# a_21080_48324# 0.00133f
C5479 AVDD a_19928_41284# 0.00159f
C5480 XA4.XA4.MN0.D a_9848_46916# 0.00396f
C5481 XA7.XA1.XA5.MN2.G a_16040_44452# 0.00486f
C5482 a_2288_48324# a_2288_47972# 0.0109f
C5483 AVDD a_14888_52900# 0.00166f
C5484 XA6.XA11.MN1.G a_11000_53604# 9.49e-20
C5485 XA5.XA11.MN1.G a_13520_53604# 0.0726f
C5486 XA5.XA1.XA1.MN0.S a_12368_39876# 2.54e-19
C5487 XA5.XA1.XA1.MN0.D a_13520_40580# 0.035f
C5488 a_2288_40932# a_2288_40580# 0.0109f
C5489 XA0.XA11.MN1.G a_13808_2798# 0.00449f
C5490 a_3440_46564# a_4808_46564# 8.89e-19
C5491 XA5.XA4.MN0.G a_13520_45156# 0.00865f
C5492 XA5.XA3.MN0.G a_13520_46564# 0.156f
C5493 a_22448_46916# a_22448_46564# 0.0109f
C5494 XA1.XA4.MN0.D a_3440_43748# 9.24e-20
C5495 AVDD a_2288_50436# 0.416f
C5496 XA1.XA10.MP0.G a_2288_52196# 0.0441f
C5497 a_7328_52548# XA3.XA9.MN1.G 0.0674f
C5498 CK_SAMPLE XA5.XA6.MN2.D 0.0389f
C5499 XA20.XA10.MN1.D XA8.XA7.MP0.G 0.00198f
C5500 XA7.XA10.MP0.G XA7.XA9.MN0.D 0.106f
C5501 XB1.XA1.MP0.D a_8408_1390# 4.8e-20
C5502 XB1.M1.G XB1.XA0.MP0.D 0.303f
C5503 XB2.XA1.MP0.D a_14960_1742# 8.72e-20
C5504 XB2.M1.G a_12368_2094# 0.00186f
C5505 SARN li_14804_28392# 0.00103f
C5506 XA7.XA4.MN0.G a_18560_42692# 0.0049f
C5507 D<1> a_17408_39876# 7.77e-20
C5508 XA20.XA3a.MN0.D XA5.XA1.XA4.MN1.D 0.0124f
C5509 XA2.XA1.XA5.MN2.D a_4808_44452# 0.153f
C5510 a_11000_45156# a_11000_44804# 0.0109f
C5511 XA20.XA2a.MN0.D a_9848_43748# 4.48e-20
C5512 a_23600_45156# XA20.XA2.MN1.D 0.00176f
C5513 XA2.XA1.XA5.MN2.G a_2288_51140# 0.0754f
C5514 AVDD a_3440_47620# 0.00125f
C5515 XA0.XA10.MP0.D VREF 0.0118f
C5516 XA2.XA9.MN1.G XA2.XA6.MP0.D 0.0618f
C5517 a_16040_51844# D<2> 1.25e-19
C5518 XA8.XA9.MN1.G a_19928_50436# 0.01f
C5519 XB1.XA4.MP0.D XDAC1.XC1.XRES1B.B 0.00184f
C5520 li_14804_25524# li_14804_24912# 0.00271f
C5521 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES2.B 0.0307f
C5522 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES16.B 0.0381f
C5523 XDAC2.XC64b<1>.XRES1A.B XDAC2.X16ab.XRES1A.B 0.00444f
C5524 XDAC1.X16ab.XRES8.B li_9184_24912# 9.91e-20
C5525 D<4> XDAC1.XC32a<0>.XRES8.B 0.00669f
C5526 XA20.XA2a.MN0.D XA8.XA1.XA1.MN0.S 0.139f
C5527 XA1.XA1.XA5.MP0.D XA1.XA1.XA5.MN0.D 0.00918f
C5528 XA5.XA1.XA5.MP1.D a_12368_43396# 0.00176f
C5529 XA1.XA1.XA2.MP0.D XA2.XA1.XA2.MP0.D 0.00435f
C5530 a_920_43748# a_920_43396# 0.0109f
C5531 EN a_920_43044# 0.141f
C5532 XA0.XA6.MP0.G XDAC2.XC128b<2>.XRES1B.B 0.00405f
C5533 XA2.XA6.MP0.G li_14804_23688# 0.00504f
C5534 a_13520_50436# a_13520_50084# 0.0109f
C5535 XA3.XA1.XA5.MN2.G a_5960_48676# 0.00363f
C5536 AVDD a_17408_44452# 0.357f
C5537 XDAC2.XC64a<0>.XRES16.B XDAC2.XC64a<0>.XRES1A.B 0.454f
C5538 EN a_n232_40580# 0.0786f
C5539 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES8.B 0.00687f
C5540 XA7.XA1.XA4.MN1.D a_18560_42340# 0.00176f
C5541 a_7328_42692# a_7328_42340# 0.0109f
C5542 D<2> a_14888_46212# 0.0141f
C5543 a_13520_49028# a_13520_48676# 0.0109f
C5544 VREF a_2288_47972# 0.0175f
C5545 D<6> a_4808_45860# 0.0675f
C5546 XA7.XA1.XA5.MN2.G a_16040_45508# 0.00595f
C5547 AVDD a_3440_41988# 0.00125f
C5548 XA5.XA4.MN0.D XA6.XA4.MN0.G 3.16e-20
C5549 XA6.XA4.MN0.D XA5.XA4.MN0.G 3.16e-20
C5550 XA20.XA12.MP0.G XA8.XA11.MN1.G 0.00369f
C5551 a_3440_53956# a_4808_53956# 8.89e-19
C5552 a_17408_54308# a_17408_53956# 0.0109f
C5553 AVDD a_920_53604# 0.383f
C5554 a_4808_54308# XA3.XA11.MN1.G 2.54e-19
C5555 XA2.XA1.XA1.MN0.S a_5960_40932# 0.0271f
C5556 a_17408_41284# a_18560_41284# 0.00133f
C5557 SARP li_9184_17952# 0.00103f
C5558 XA5.XA1.XA5.MN2.G XA5.XA1.XA4.MP1.D 7.44e-19
C5559 D<7> a_2288_43044# 7.77e-20
C5560 a_8480_47268# a_8480_46916# 0.0109f
C5561 VREF a_16040_44804# 0.0691f
C5562 AVDD a_9560_2094# 0.00154f
C5563 D<3> a_12368_43396# 7.77e-20
C5564 XA1.XA6.MP0.G a_2288_43748# 5.5e-19
C5565 AVDD XA8.XA1.XA5.MN2.G 4.81f
C5566 XA0.XA10.MP0.D a_920_52548# 0.00224f
C5567 a_12368_52900# a_13520_52900# 0.00133f
C5568 a_920_52900# XA0.XA10.MP0.G 0.0658f
C5569 CK_SAMPLE XA3.XA8.MP0.D 3.93e-19
C5570 XA0.XA12.MP0.D a_2288_51844# 4.48e-19
C5571 DONE a_21080_51492# 0.00837f
C5572 a_8408_3502# a_9560_3502# 0.00133f
C5573 XA20.XA3a.MN0.D XA2.XA1.XA5.MN0.D 0.0106f
C5574 a_4808_45508# XA2.XA1.XA5.MN2.D 0.0674f
C5575 XA3.XA4.MN0.G a_7328_43396# 8.07e-19
C5576 XA5.XA1.XA5.MN2.G a_11000_40228# 0.0108f
C5577 XA8.XA3.MN0.G a_21080_44452# 0.055f
C5578 XA1.XA3.MN0.G a_4808_44100# 4.4e-20
C5579 XA2.XA3.MN0.G a_3440_44100# 4.21e-19
C5580 AVDD a_2288_48676# 0.356f
C5581 CK_SAMPLE a_12368_49380# 7.89e-19
C5582 XA7.XA9.MN1.G a_17408_51140# 0.0222f
C5583 a_22448_51844# a_23600_51844# 0.00133f
C5584 XA6.XA7.MP0.D a_14888_51492# 0.124f
C5585 a_22448_53956# VREF 0.0012f
C5586 D<5> XDAC1.X16ab.XRES2.B 0.00405f
C5587 EN XA7.XA1.XA5.MN1.D 0.0157f
C5588 XA7.XA1.XA5.MN2.D a_17408_43044# 1.88e-19
C5589 XA20.XA2a.MN0.D a_5960_42340# 0.00732f
C5590 a_5960_51492# VREF 0.00396f
C5591 a_920_50788# XA0.XA6.MP0.G 1.34e-19
C5592 a_n232_50436# a_920_50436# 0.00133f
C5593 AVDD a_17408_45508# 0.359f
C5594 XA1.XA1.XA2.MP0.D a_3440_41988# 0.0568f
C5595 XA5.XA1.XA2.MP0.D a_13520_42340# 0.0966f
C5596 a_11000_43044# a_11000_42692# 0.0109f
C5597 XA1.XA4.MN0.D XDAC1.XC32a<0>.XRES1A.A 0.0216f
C5598 XA4.XA1.XA5.MN2.G a_7328_46564# 0.00363f
C5599 a_5960_49380# a_7328_49380# 8.89e-19
C5600 XA3.XA6.MP0.G XA3.XA4.MN0.G 0.0407f
C5601 AVDD XA4.XA1.XA4.MP1.D 0.0913f
C5602 XA0.XA4.MN0.D a_920_49028# 0.154f
C5603 VREF a_n232_49028# 7.81e-19
C5604 AVDD a_23600_55364# 0.00236f
C5605 a_14888_47972# a_14888_47620# 0.0109f
C5606 XA4.XA4.MN0.G a_11000_47268# 0.155f
C5607 a_920_47620# a_2288_47620# 8.89e-19
C5608 XA0.XA6.MP2.G a_920_43748# 7.76e-20
C5609 XA3.XA1.XA5.MN2.G XA2.XA1.XA5.MP0.D 0.00353f
C5610 XA4.XA4.MN0.D a_9848_45860# 5.88e-20
C5611 XA7.XA6.MP0.G a_17408_45156# 5.5e-19
C5612 VREF a_14888_45860# 1.19e-19
C5613 AVDD a_9848_40228# 0.00131f
C5614 XA7.XA12.MP0.G a_17408_52900# 1.28e-19
C5615 XA8.XA11.MN1.G a_18560_52900# 0.00295f
C5616 XA6.XA11.MP0.D a_16040_53252# 0.0494f
C5617 CK_SAMPLE XA0.XA9.MN1.G 0.134f
C5618 AVDD a_16040_52196# 0.37f
C5619 XA4.XA11.MN1.G XA3.XA10.MP0.G 0.00598f
C5620 XA0.XA11.MN1.G XA0.XA10.MP0.D 0.0625f
C5621 a_21080_40580# a_21080_40228# 0.0109f
C5622 XA20.XA3a.MN0.D a_18560_44452# 2.59e-20
C5623 XA8.XA3.MN0.G a_21080_45508# 0.0698f
C5624 XA0.XA7.MP0.G XA0.XA1.XA1.MN0.D 0.0384f
C5625 XA7.XA1.XA5.MN2.G a_17408_41284# 5.96e-19
C5626 XA4.XA6.MP0.G XA4.XA1.XA4.MP0.D 9.97e-19
C5627 XA2.XA4.MN0.D a_5960_43044# 9.14e-20
C5628 XA4.XA4.MN0.G EN 0.0579f
C5629 XA8.XA4.MN0.G a_19928_44100# 0.0164f
C5630 XA1.XA4.MN0.G XA1.XA1.XA5.MP1.D 0.00138f
C5631 a_21080_46212# a_22448_46212# 8.89e-19
C5632 XA5.XA10.MP0.G a_13520_51492# 6.8e-20
C5633 AVDD a_920_49732# 0.359f
C5634 CK_SAMPLE XA6.XA6.MP0.D 0.0276f
C5635 XA3.XA9.MN0.D a_8480_51844# 0.00176f
C5636 XA3.XA9.MN1.G a_9848_51844# 2.2e-19
C5637 a_3440_52196# XA1.XA7.MP0.D 0.0662f
C5638 XA8.XA9.MN1.G XA7.XA7.MP0.D 0.00108f
C5639 a_13808_686# CK_SAMPLE_BSSW 0.0709f
C5640 XB2.XA3.MN1.D m3_26048_132# 0.17f
C5641 a_14888_44452# a_16040_44452# 0.00133f
C5642 SARN XDAC2.XC128a<1>.XRES8.B 27.7f
C5643 XA20.XA3a.MN0.D a_4808_41988# 0.00547f
C5644 XA20.XA2a.MN0.D a_13520_43044# 1.43e-19
C5645 a_7328_44804# EN 3.4e-19
C5646 XA2.XA4.MN0.D a_4808_40580# 9.25e-20
C5647 XA5.XA9.MN1.G VREF 0.0732f
C5648 AVDD a_4808_46564# 0.00125f
C5649 XA8.XA7.MP0.G a_22448_50788# 0.0012f
C5650 D<5> D<3> 0.00362f
C5651 D<7> D<1> 4.29e-19
C5652 XA0.XA9.MN1.G a_920_49380# 2.54e-19
C5653 D<6> D<2> 0.184f
C5654 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128a<1>.XRES8.B 6.7e-19
C5655 XB2.XA3.MN1.D m3_16472_3476# 0.0137f
C5656 li_9184_20208# li_9184_19596# 0.00271f
C5657 XA0.XA4.MN0.D XDAC1.XC128b<2>.XRES1B.B 0.00405f
C5658 XA4.XA6.MP0.G li_14804_14472# 0.00504f
C5659 XA0.XA6.MP0.G li_14804_12636# 1.76e-19
C5660 EN XA6.XA1.XA4.MP0.D 0.0386f
C5661 a_14888_43396# a_16040_43396# 0.00133f
C5662 XA0.XA6.MP0.G a_920_49028# 0.0307f
C5663 XA8.XA7.MP0.G XA20.XA3a.MN0.D 0.203f
C5664 D<6> XA2.XA4.MN0.G 0.259f
C5665 XA3.XA1.XA5.MN2.G a_5960_47620# 0.00363f
C5666 AVDD XA1.XA1.XA5.MN0.D 0.00889f
C5667 XA4.XA6.MP0.G a_11000_49380# 0.0781f
C5668 a_920_41988# a_2288_41988# 8.89e-19
C5669 D<6> a_4808_44804# 5.24e-19
C5670 a_9848_48324# XA4.XA4.MN0.G 0.0677f
C5671 AVDD a_18560_41284# 0.00125f
C5672 XA7.XA1.XA5.MN2.G a_14888_44452# 1.86e-19
C5673 D<2> a_16040_45156# 6.68e-19
C5674 AVDD a_13520_52900# 0.00166f
C5675 a_23600_53956# a_23600_53604# 0.0109f
C5676 XA4.XA12.MP0.G a_11000_53604# 0.0893f
C5677 XA5.XA11.MN1.G a_12368_53604# 0.073f
C5678 SARP XDAC1.XC1.XRES8.B 27.7f
C5679 XA5.XA1.XA1.MN0.D a_12368_40580# 8.3e-19
C5680 a_13520_40932# a_14888_40932# 8.89e-19
C5681 XA0.XA11.MN1.G a_12368_2798# 0.0947f
C5682 XA5.XA4.MN0.G a_12368_45156# 5.54e-19
C5683 XA5.XA3.MN0.G a_12368_46564# 0.155f
C5684 XA3.XA1.XA5.MN2.G a_5960_41988# 0.0719f
C5685 XA1.XA4.MN0.D a_2288_43748# 9.15e-20
C5686 AVDD a_920_50436# 0.416f
C5687 CK_SAMPLE XA5.XA6.MP2.D 3.06e-19
C5688 a_18560_52548# a_19928_52548# 8.89e-19
C5689 XA7.XA10.MP0.G XA7.XA9.MN1.G 0.202f
C5690 SAR_IP XB1.XA3.MN1.D 0.234f
C5691 SAR_IN a_14960_1742# 0.0215f
C5692 XB2.XA1.MP0.D a_13808_1742# 8.33e-19
C5693 XA4.XA3.MN0.G XA4.XA1.XA2.MP0.D 0.00212f
C5694 XA7.XA4.MN0.G a_17408_42692# 0.00224f
C5695 XA20.XA3a.MN0.D XA5.XA1.XA4.MP1.D 0.0124f
C5696 XA20.XA2a.MN0.D a_8480_43748# 2.91e-20
C5697 XA0.XA7.MP0.G a_2288_51140# 7.1e-20
C5698 XA2.XA1.XA5.MN2.G a_920_51140# 7.1e-20
C5699 a_13520_51492# a_13520_51140# 0.0109f
C5700 AVDD a_2288_47620# 0.356f
C5701 XA6.XA1.XA5.MN2.G XA7.XA1.XA5.MN2.G 0.0255f
C5702 XA4.XA7.MP0.D a_9848_50788# 3.29e-19
C5703 XA2.XA9.MN1.G XA2.XA6.MN0.D 0.0615f
C5704 XA20.XA2a.MN0.D XA7.XA1.XA1.MP2.D 0.0102f
C5705 XA1.XA1.XA2.MP0.D XA1.XA1.XA5.MN0.D 0.056f
C5706 a_13520_43748# XA5.XA1.XA5.MN0.D 0.00176f
C5707 D<3> XDAC1.XC32a<0>.XRES4.B 0.00405f
C5708 XA2.XA3.MN0.G XA2.XA1.XA1.MN0.D 0.00135f
C5709 EN a_n232_43044# 0.0754f
C5710 XA0.XA6.MN0.D a_n232_50084# 0.0488f
C5711 XA0.XA6.MP0.G a_920_50084# 0.159f
C5712 XA8.XA7.MP0.G a_22448_49028# 8.22e-19
C5713 XA5.XA6.MP0.G XA5.XA6.MP0.D 0.0392f
C5714 XA8.XA6.MP2.D VREF 6.11e-19
C5715 AVDD a_16040_44452# 0.357f
C5716 D<8> XDAC2.XC64b<1>.XRES8.B 4.06e-21
C5717 a_18560_42692# XA7.XA1.XA4.MN0.D 0.00176f
C5718 a_n232_48676# a_920_48676# 0.00133f
C5719 VREF a_920_47972# 0.0175f
C5720 D<6> a_3440_45860# 1.06e-19
C5721 XA7.XA1.XA5.MN2.G a_14888_45508# 2.31e-19
C5722 AVDD a_2288_41988# 0.386f
C5723 XA5.XA4.MN0.D XA5.XA4.MN0.G 0.707f
C5724 AVDD a_n232_53604# 0.00166f
C5725 a_23600_55364# XA20.XA10.MN1.D 8.48e-20
C5726 XA6.XA1.XA1.MP2.D XA6.XA1.XA1.MP1.D 0.0488f
C5727 a_4808_41284# XA2.XA1.XA1.MN0.D 0.00224f
C5728 AVDD a_8408_2094# 0.362f
C5729 XA4.XA4.MN0.G a_11000_46212# 3.46e-19
C5730 XA5.XA1.XA5.MN2.G XA4.XA1.XA4.MP1.D 0.00353f
C5731 a_19928_47268# a_21080_47268# 0.00133f
C5732 VREF a_14888_44804# 7.12e-19
C5733 AVDD XA7.XA1.XA5.MN2.G 5.46f
C5734 a_n232_53252# XA0.XA9.MN1.G 5.25e-19
C5735 XA0.XA10.MP0.D a_n232_52548# 0.00316f
C5736 a_n232_52900# XA0.XA10.MP0.G 0.0681f
C5737 XA5.XA10.MP0.D XA5.XA10.MP0.G 0.194f
C5738 CK_SAMPLE XA2.XA8.MP0.D 3.93e-19
C5739 XA0.XA12.MP0.D a_920_51844# 2.62e-19
C5740 DONE a_19928_51492# 0.00357f
C5741 a_9560_3854# a_9560_3502# 0.0109f
C5742 XA20.XA3a.MN0.D XA2.XA1.XA2.MP0.D 0.195f
C5743 a_21080_45860# XA8.XA1.XA5.MN2.D 3.12e-20
C5744 a_14888_45508# a_16040_45508# 0.00133f
C5745 XA5.XA1.XA5.MN2.G a_9848_40228# 5.59e-19
C5746 SARN a_13808_1742# 9.76e-19
C5747 XA0.XA4.MN0.D a_920_42340# 9.14e-20
C5748 XA1.XA3.MN0.G a_3440_44100# 0.00776f
C5749 XA8.XA3.MN0.G a_19928_44452# 0.0934f
C5750 AVDD a_920_48676# 0.356f
C5751 XA1.XA9.MN1.G XA1.XA6.MN2.D 0.126f
C5752 CK_SAMPLE a_11000_49380# 7.89e-19
C5753 a_4808_51844# a_4808_51492# 0.0109f
C5754 a_13520_51844# XA5.XA8.MP0.D 0.0215f
C5755 a_21080_53956# VREF 0.00311f
C5756 li_14804_30648# li_14804_30036# 0.00271f
C5757 XDAC2.XC0.XRES8.B XDAC2.XC64b<1>.XRES8.B 6.7e-19
C5758 SARN li_14804_8124# 0.00103f
C5759 a_9848_44100# a_9848_43748# 0.0109f
C5760 a_21080_44100# XA8.XA1.XA5.MP1.D 0.00176f
C5761 EN XA7.XA1.XA5.MP1.D 0.0543f
C5762 XA20.XA3a.MN0.D a_19928_41284# 0.00649f
C5763 XA20.XA2a.MN0.D a_4808_42340# 0.0843f
C5764 a_8480_44452# XA3.XA1.XA2.MP0.D 5.16e-20
C5765 XA3.XA1.XA5.MP1.D XA3.XA1.XA5.MN1.D 0.00918f
C5766 XA0.XA6.MP2.G XDAC1.X16ab.XRES1A.B 4.06e-21
C5767 XA8.XA7.MP0.G a_22448_50084# 0.00104f
C5768 D<2> XA3.XA6.MP0.G 0.0286f
C5769 a_n232_50788# XA0.XA6.MP0.G 1.75e-20
C5770 a_12368_50788# a_12368_50436# 0.0109f
C5771 D<4> XA5.XA6.MP0.G 9.98e-20
C5772 D<1> XA2.XA6.MP0.G 0.037f
C5773 D<3> XA4.XA6.MP0.G 0.0523f
C5774 AVDD a_16040_45508# 0.359f
C5775 XDAC2.XC32a<0>.XRES4.B XDAC2.XC32a<0>.XRES8.B 0.471f
C5776 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES2.B 0.0136f
C5777 XA5.XA1.XA2.MP0.D a_12368_42340# 2.54e-19
C5778 XA1.XA1.XA2.MP0.D a_2288_41988# 0.0219f
C5779 EN XA2.XA1.XA1.MN0.S 0.139f
C5780 XA6.XA6.MP0.G a_16040_48324# 0.00417f
C5781 XA4.XA1.XA5.MN2.G a_5960_46564# 7.1e-20
C5782 XA3.XA1.XA5.MN2.G a_7328_46564# 7.1e-20
C5783 AVDD XA4.XA1.XA4.MN1.D 0.00889f
C5784 XA0.XA4.MN0.D a_n232_49028# 0.156f
C5785 XA6.XA4.MN0.D a_16040_49380# 0.154f
C5786 AVDD a_22448_55364# 0.448f
C5787 SARP li_9184_28392# 0.00103f
C5788 a_21080_41988# XA8.XA1.XA1.MN0.S 3.8e-19
C5789 a_19928_41636# a_21080_41636# 0.00133f
C5790 a_8480_41636# XA3.XA1.XA1.MN0.S 0.0658f
C5791 a_7328_41636# XA3.XA1.XA1.MP2.D 0.00176f
C5792 XA4.XA4.MN0.G a_9848_47268# 0.157f
C5793 XA0.XA6.MP2.G a_n232_43748# 6.49e-19
C5794 XA3.XA1.XA5.MN2.G XA2.XA1.XA5.MN0.D 7.2e-19
C5795 VREF a_13520_45860# 1.19e-19
C5796 AVDD a_8480_40228# 0.00131f
C5797 AVDD a_14888_52196# 0.00154f
C5798 XA8.XA11.MN1.G a_17408_52900# 1.34e-19
C5799 a_4808_53252# a_5960_53252# 0.00133f
C5800 CK_SAMPLE a_23600_52548# 8.45e-19
C5801 a_7328_40228# a_8480_40228# 0.00133f
C5802 XA2.XA3.MN0.G XA2.XA1.XA5.MN2.D 0.753f
C5803 XA8.XA3.MN0.G a_19928_45508# 0.104f
C5804 XA4.XA6.MP0.G XA4.XA1.XA4.MN0.D 6.07e-19
C5805 XA7.XA1.XA5.MN2.G a_16040_41284# 0.0175f
C5806 XA2.XA4.MN0.D a_4808_43044# 9.25e-20
C5807 XA3.XA4.MN0.G EN 0.0578f
C5808 XA7.XA4.MN0.G a_19928_44100# 2.84e-19
C5809 XA8.XA4.MN0.G a_18560_44100# 2.84e-19
C5810 XA0.XA6.MP0.G a_920_42340# 5.5e-19
C5811 SARN a_23600_40228# 9.45e-19
C5812 a_8480_46212# a_8480_45860# 0.0109f
C5813 a_12368_52900# XA6.XA1.XA5.MN2.G 1.06e-19
C5814 CK_SAMPLE XA6.XA6.MN0.D 0.0659f
C5815 XA7.XA9.MN1.G XA8.XA7.MP0.D 0.00108f
C5816 XA7.XA9.MN0.D XA7.XA7.MP0.D 0.00986f
C5817 AVDD a_n232_49732# 0.00159f
C5818 XA3.XA9.MN1.G a_8480_51844# 0.0164f
C5819 a_2288_52196# XA1.XA7.MP0.D 0.0674f
C5820 a_13520_52196# a_14888_52196# 8.89e-19
C5821 a_13808_686# a_14960_686# 0.00133f
C5822 a_9560_686# a_9560_334# 0.0109f
C5823 XB2.XA3.MN1.D m3_25976_132# 0.0634f
C5824 XA20.XA3a.MN0.D a_3440_41988# 0.00547f
C5825 XA5.XA1.XA5.MN2.D a_13520_43748# 0.00224f
C5826 XA4.XA4.MN0.G a_9848_41636# 6.69e-20
C5827 a_2288_44452# a_2288_44100# 0.0109f
C5828 a_5960_44804# EN 3.4e-19
C5829 XA3.XA9.MN1.G XA3.XA4.MN0.D 0.00938f
C5830 a_2288_51492# XA1.XA6.MP0.G 4.06e-20
C5831 AVDD a_3440_46564# 0.00125f
C5832 XA8.XA7.MP0.G a_21080_50788# 0.00548f
C5833 a_9848_51140# a_9848_50788# 0.0109f
C5834 a_21080_51140# XA8.XA6.MP2.D 0.00176f
C5835 XA0.XA9.MN1.G a_n232_49380# 4.23e-20
C5836 XA4.XA7.MP0.D a_9848_50084# 7.44e-20
C5837 XB2.XA3.MN1.D m3_26048_4356# 0.17f
C5838 XA0.XA6.MP0.G XDAC2.XC32a<0>.XRES1A.A 0.00169f
C5839 EN XA6.XA1.XA4.MN0.D 3.17e-19
C5840 XA7.XA6.MP0.G XDAC2.XC32a<0>.XRES1B.B 0.00405f
C5841 XA5.XA6.MP0.G li_14804_15084# 0.00504f
C5842 XA6.XA1.XA2.MP0.D a_16040_43044# 3.59e-19
C5843 XA2.XA1.XA2.MP0.D XA2.XA1.XA4.MP1.D 4.34e-19
C5844 XA6.XA1.XA5.MN0.D a_14888_43044# 0.00176f
C5845 a_2288_43396# a_2288_43044# 0.0109f
C5846 a_12368_50084# a_12368_49732# 0.0109f
C5847 a_n232_50084# XA0.XA4.MN0.D 3.12e-20
C5848 XA0.XA6.MP0.G a_n232_49028# 0.0137f
C5849 XA8.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.96f
C5850 XA20.XA3.MN1.D VREF 0.00124f
C5851 AVDD XA1.XA1.XA5.MP0.D 0.159f
C5852 XA4.XA6.MP0.G a_9848_49380# 0.0547f
C5853 SARP a_13808_1742# 2.97e-20
C5854 D<8> li_14804_18564# 0.00508f
C5855 a_13520_42340# a_13520_41988# 0.0109f
C5856 a_18560_48324# a_19928_48324# 8.89e-19
C5857 AVDD a_17408_41284# 0.361f
C5858 VREF a_12368_46916# 0.0536f
C5859 XA3.XA4.MN0.D a_8480_46916# 0.00456f
C5860 XA6.XA1.XA5.MN2.G a_14888_44452# 5.11e-19
C5861 D<2> a_14888_45156# 7.77e-19
C5862 a_920_48324# a_920_47972# 0.0109f
C5863 AVDD a_12368_52900# 0.387f
C5864 XA4.XA12.MP0.G a_9848_53604# 0.1f
C5865 XA5.XA11.MN1.G a_11000_53604# 0.0124f
C5866 XA0.XA1.XA1.MN0.D a_n232_40228# 0.00155f
C5867 XA5.XA1.XA1.MP1.D a_12368_40580# 0.00176f
C5868 a_920_40932# a_920_40580# 0.0109f
C5869 XA0.XA11.MN1.G a_11000_2798# 0.0931f
C5870 D<5> XA3.XA1.XA4.MN0.D 0.00144f
C5871 a_2288_46564# a_3440_46564# 0.00133f
C5872 a_21080_46916# a_21080_46564# 0.0109f
C5873 XA8.XA7.MP0.G a_22448_42340# 9.75e-19
C5874 XA3.XA1.XA5.MN2.G a_4808_41988# 0.0684f
C5875 D<1> a_18560_42692# 6.49e-19
C5876 VREF a_2288_43748# 8.43e-19
C5877 CK_SAMPLE D<3> 0.0524f
C5878 AVDD a_n232_50436# 0.00154f
C5879 XA0.XA10.MP0.G a_920_52196# 0.0441f
C5880 XB1.XA1.MN0.D XB1.XA3.MN1.D 2.08e-19
C5881 a_14960_2798# XB2.XA3.MN1.D 3.55e-19
C5882 a_14960_2446# a_14960_2094# 0.0109f
C5883 SAR_IP XB1.XA3.MN0.S 0.0903f
C5884 SAR_IN a_13808_1742# 0.0425f
C5885 SARN XDAC2.XC64b<1>.XRES8.B 27.7f
C5886 XA3.XA3.MN0.G XA4.XA1.XA2.MP0.D 0.00485f
C5887 XA0.XA4.MN0.G XA0.XA1.XA4.MN0.D 0.00331f
C5888 XA5.XA6.MP0.G a_13520_40932# 3.97e-20
C5889 XA20.XA3a.MN0.D XA4.XA1.XA4.MP1.D 0.0124f
C5890 XA1.XA1.XA5.MN2.D a_3440_44452# 0.153f
C5891 XA8.XA1.XA5.MN2.D a_21080_44804# 0.156f
C5892 a_9848_45156# a_9848_44804# 0.0109f
C5893 a_22448_45156# a_23600_45156# 0.00133f
C5894 XA1.XA6.MP0.G a_3440_40580# 7.76e-20
C5895 a_920_51492# XA0.XA6.MP2.G 2.41e-19
C5896 XA0.XA7.MP0.G a_920_51140# 0.077f
C5897 AVDD a_920_47620# 0.356f
C5898 a_22448_53252# VREF 0.00125f
C5899 XA2.XA9.MN1.G XA2.XA6.MP0.G 0.0725f
C5900 li_9184_25524# li_9184_24912# 0.00271f
C5901 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES2.B 0.0307f
C5902 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES16.B 0.0381f
C5903 XDAC1.XC64b<1>.XRES1A.B XDAC1.X16ab.XRES1A.B 0.00444f
C5904 XA20.XA2a.MN0.D XA7.XA1.XA1.MN0.S 0.137f
C5905 XA1.XA1.XA2.MP0.D XA1.XA1.XA5.MP0.D 4.34e-19
C5906 XA4.XA1.XA5.MP1.D a_11000_43396# 0.00176f
C5907 a_n232_43748# a_n232_43396# 0.0109f
C5908 XA2.XA6.MP0.G XDAC2.X16ab.XRES16.B 0.0181f
C5909 a_12368_50436# a_12368_50084# 0.0109f
C5910 XA0.XA6.MP0.G a_n232_50084# 6.4e-20
C5911 XA8.XA7.MP0.G a_21080_49028# 0.00363f
C5912 XA4.XA6.MP0.G XA6.XA6.MP0.G 0.321f
C5913 XA3.XA6.MP0.G XA7.XA6.MP0.G 0.0316f
C5914 D<5> a_8480_49380# 5.91e-19
C5915 AVDD a_14888_44452# 0.00125f
C5916 XDAC1.XC64a<0>.XRES16.B XDAC1.XC64a<0>.XRES1A.B 0.454f
C5917 XDAC2.XC64a<0>.XRES16.B li_14804_9768# 0.00117f
C5918 XA1.XA3.MN0.G li_14804_29004# 0.00504f
C5919 EN a_22448_40932# 5.7e-20
C5920 SARP a_23600_40228# 0.0038f
C5921 XA7.XA1.XA2.MP0.D XA7.XA1.XA1.MN0.S 2.11e-19
C5922 XA2.XA1.XA4.MN0.D XA2.XA1.XA4.MP0.D 0.00918f
C5923 XA7.XA1.XA4.MP1.D a_17408_42340# 0.00176f
C5924 a_5960_42692# a_5960_42340# 0.0109f
C5925 XA2.XA6.MP0.G a_5960_46916# 5.5e-19
C5926 XA6.XA6.MP0.G a_16040_47268# 5.95e-19
C5927 a_12368_49028# a_12368_48676# 0.0109f
C5928 XA0.XA4.MN0.D a_920_47972# 0.0546f
C5929 XA6.XA1.XA5.MN2.G a_14888_45508# 9.01e-20
C5930 AVDD a_920_41988# 0.386f
C5931 VREF a_n232_47972# 7.39e-19
C5932 a_4808_54308# XA2.XA11.MN1.G 2.9e-19
C5933 AVDD XA20.XA10.MN0.D 4.25e-19
C5934 a_16040_54308# a_16040_53956# 0.0109f
C5935 a_2288_53956# a_3440_53956# 0.00133f
C5936 XA6.XA1.XA1.MN0.S XA6.XA1.XA1.MP1.D 0.0615f
C5937 a_16040_41284# a_17408_41284# 8.89e-19
C5938 SARP XDAC1.XC128a<1>.XRES8.B 27.7f
C5939 AVDD XB2.XA4.MP0.D 2.39f
C5940 VREF a_13520_44804# 7.12e-19
C5941 XA4.XA6.MP0.G XA4.XA1.XA5.MP1.D 0.00121f
C5942 XA5.XA1.XA5.MN2.G XA4.XA1.XA4.MN1.D 7.2e-19
C5943 XA4.XA1.XA5.MN2.G XA4.XA1.XA4.MP1.D 7.44e-19
C5944 a_7328_47268# a_7328_46916# 0.0109f
C5945 XA4.XA4.MN0.G a_9848_46212# 0.0149f
C5946 CK_SAMPLE XA1.XA8.MP0.D 3.93e-19
C5947 AVDD XA6.XA1.XA5.MN2.G 4.81f
C5948 XA8.XA11.MN1.G a_18560_52196# 1.84e-19
C5949 a_11000_52900# a_12368_52900# 8.89e-19
C5950 XA4.XA11.MN1.G XA3.XA7.MP0.D 4.87e-19
C5951 XA20.XA3a.MN0.D XA1.XA1.XA5.MN0.D 0.0107f
C5952 a_3440_45508# XA1.XA1.XA5.MN2.D 0.0658f
C5953 XA6.XA6.MP0.G a_16040_41636# 5.5e-19
C5954 XA2.XA4.MN0.G a_5960_43396# 8.07e-19
C5955 XA8.XA4.MN0.G XA8.XA1.XA5.MP0.D 0.00138f
C5956 XA4.XA1.XA5.MN2.G a_9848_40228# 0.0709f
C5957 SARN a_12368_1742# 0.00741f
C5958 XA0.XA4.MN0.D a_n232_42340# 9.25e-20
C5959 XA1.XA3.MN0.G a_2288_44100# 0.00245f
C5960 AVDD a_n232_48676# 0.00129f
C5961 XA1.XA9.MN1.G XA1.XA6.MP2.D 0.0618f
C5962 CK_SAMPLE a_9848_49380# 0.00139f
C5963 a_12368_51844# XA5.XA8.MP0.D 0.0215f
C5964 a_21080_51844# a_22448_51844# 8.89e-19
C5965 XA5.XA7.MP0.D a_13520_51492# 0.126f
C5966 EN XA6.XA1.XA5.MP1.D 0.0544f
C5967 XA20.XA3a.MN0.D a_18560_41284# 0.00649f
C5968 XA6.XA1.XA5.MN2.D a_16040_43044# 1.88e-19
C5969 XA20.XA2a.MN0.D a_3440_42340# 0.0848f
C5970 a_18560_44804# XA7.XA1.XA2.MP0.D 2.6e-20
C5971 XA8.XA7.MP0.G a_21080_50084# 0.00366f
C5972 D<4> XA4.XA6.MP0.D 0.0323f
C5973 AVDD a_14888_45508# 0.00131f
C5974 a_21080_43044# XA8.XA1.XA4.MP1.D 0.00176f
C5975 a_9848_43044# a_9848_42692# 0.0109f
C5976 XA0.XA4.MN0.D XDAC1.XC32a<0>.XRES1A.A 0.00169f
C5977 XA6.XA6.MP0.G a_14888_48324# 0.00295f
C5978 XA8.XA7.MP0.G XA8.XA3.MN0.G 0.106f
C5979 XA3.XA1.XA5.MN2.G a_5960_46564# 0.00363f
C5980 a_4808_49380# a_5960_49380# 0.00133f
C5981 XA0.XA6.MP0.G a_920_47972# 8.92e-19
C5982 AVDD XA3.XA1.XA4.MN1.D 0.00889f
C5983 VREF a_22448_49380# 0.00186f
C5984 XA6.XA4.MN0.D a_14888_49380# 0.155f
C5985 a_7328_41636# XA3.XA1.XA1.MN0.S 0.071f
C5986 a_13520_47972# a_13520_47620# 0.0109f
C5987 a_n232_47620# a_920_47620# 0.00133f
C5988 D<2> EN 0.0683f
C5989 XA3.XA1.XA5.MN2.G XA2.XA1.XA2.MP0.D 0.144f
C5990 VREF a_12368_45860# 0.0178f
C5991 XA3.XA4.MN0.D a_8480_45860# 2.23e-19
C5992 AVDD a_7328_40228# 0.464f
C5993 AVDD a_13520_52196# 0.00154f
C5994 XA7.XA11.MN1.G a_18560_52900# 0.00208f
C5995 CK_SAMPLE a_22448_52548# 0.00672f
C5996 XA3.XA11.MN1.G XA3.XA10.MP0.G 0.0119f
C5997 a_14888_53604# XA6.XA10.MP0.D 1.17e-19
C5998 a_23600_53604# a_23600_53252# 0.0109f
C5999 a_19928_40580# a_19928_40228# 0.0109f
C6000 XA2.XA3.MN0.G XA1.XA1.XA5.MN2.D 0.00786f
C6001 XA1.XA3.MN0.G XA2.XA1.XA5.MN2.D 4.26e-19
C6002 XA0.XA4.MN0.G XA0.XA1.XA5.MP1.D 0.00138f
C6003 XA7.XA4.MN0.G a_18560_44100# 0.0164f
C6004 XA2.XA4.MN0.G EN 0.0579f
C6005 XA7.XA1.XA5.MN2.G a_14888_41284# 0.00527f
C6006 XA0.XA6.MP0.G a_n232_42340# 7.76e-20
C6007 a_19928_46212# a_21080_46212# 0.00133f
C6008 CK_SAMPLE XA6.XA6.MP0.G 0.046f
C6009 XA7.XA9.MN1.G XA7.XA7.MP0.D 0.274f
C6010 AVDD XA20.XA3.MN0.D 0.628f
C6011 XA3.XA9.MN1.G a_7328_51844# 6.57e-19
C6012 XA5.XA1.XA5.MN2.D a_12368_43748# 0.00388f
C6013 D<8> a_n232_42692# 0.00335f
C6014 a_13520_44452# a_14888_44452# 8.89e-19
C6015 a_4808_44804# EN 7.78e-19
C6016 XA7.XA6.MP0.G a_18560_39876# 7.76e-20
C6017 XA1.XA4.MN0.D a_3440_40580# 9.24e-20
C6018 SARN li_14804_18564# 0.00103f
C6019 XA4.XA9.MN1.G VREF 0.0732f
C6020 AVDD a_2288_46564# 0.356f
C6021 XA8.XA7.MP0.G a_19928_50788# 1.87e-19
C6022 XA7.XA9.MN1.G a_18560_49732# 0.00119f
C6023 XB2.XA3.MN1.D m3_25976_4356# 0.0634f
C6024 XDAC2.XC128b<2>.XRES16.B XDAC2.XC128b<2>.XRES1A.B 0.454f
C6025 XA4.XA6.MP0.G XDAC2.XC32a<0>.XRES8.B 0.00669f
C6026 EN XA5.XA1.XA4.MN0.D 3.17e-19
C6027 XA20.XA2a.MN0.D a_9848_40580# 0.00138f
C6028 XA2.XA1.XA2.MP0.D XA2.XA1.XA4.MN1.D 0.056f
C6029 XA6.XA1.XA2.MP0.D a_14888_43044# 0.0292f
C6030 a_13520_43396# a_14888_43396# 8.89e-19
C6031 XA7.XA6.MP0.G XA7.XA4.MN0.D 0.76f
C6032 XA8.XA7.MP0.G a_22448_47972# 8.22e-19
C6033 XA7.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.885f
C6034 D<3> a_13520_48324# 6.53e-19
C6035 XA20.XA3.MN6.D VREF 0.0398f
C6036 AVDD XA1.XA1.XA2.MP0.D 0.263f
C6037 SARP a_12368_1742# 0.0369f
C6038 a_12368_42692# XA5.XA1.XA1.MN0.S 6.76e-20
C6039 a_n232_41988# a_920_41988# 0.00133f
C6040 a_8480_48324# XA3.XA4.MN0.G 0.0661f
C6041 XA6.XA1.XA5.MN2.G a_13520_44452# 1.86e-19
C6042 AVDD a_16040_41284# 0.361f
C6043 VREF a_11000_46916# 0.0536f
C6044 XA3.XA4.MN0.D a_7328_46916# 0.00254f
C6045 XA2.XA6.MP0.G a_5960_45860# 5.5e-19
C6046 XA6.XA6.MP0.G a_16040_46212# 5.5e-19
C6047 XA20.XA10.MN1.D XA20.XA10.MN0.D 0.142f
C6048 AVDD a_11000_52900# 0.387f
C6049 DONE XA20.XA9.MP0.D 0.00306f
C6050 a_22448_53956# a_22448_53604# 0.0109f
C6051 XA5.XA11.MN1.G a_9848_53604# 0.00305f
C6052 SARP li_9184_8124# 0.00103f
C6053 XA4.XA1.XA1.MN0.S a_11000_39876# 2.54e-19
C6054 a_12368_40932# a_13520_40932# 0.00133f
C6055 XA0.XA11.MN1.G a_9560_2798# 0.00449f
C6056 D<5> XA3.XA1.XA4.MP0.D 6.09e-19
C6057 XA5.XA6.MP0.G a_13520_43396# 7.76e-20
C6058 XA1.XA6.MP0.G a_3440_43044# 7.76e-20
C6059 XA4.XA4.MN0.G a_11000_45156# 5.54e-19
C6060 XA4.XA3.MN0.G a_11000_46564# 0.155f
C6061 XA8.XA7.MP0.G a_21080_42340# 0.00442f
C6062 D<1> a_17408_42692# 7.77e-20
C6063 XA2.XA1.XA5.MN2.G a_4808_41988# 0.00407f
C6064 VREF a_920_43748# 8.43e-19
C6065 a_17408_52548# a_18560_52548# 0.00133f
C6066 XA6.XA10.MP0.G XA6.XA9.MN0.D 0.106f
C6067 AVDD a_23600_50788# 0.00181f
C6068 CK_SAMPLE XA4.XA6.MP2.D 3.06e-19
C6069 a_4808_52548# XA2.XA9.MN0.D 0.00176f
C6070 a_5960_52548# XA2.XA9.MN1.G 0.0658f
C6071 XA0.XA10.MP0.G a_n232_52196# 0.0131f
C6072 XB1.XA1.MP0.D XB1.XA3.MN1.D 4.9e-19
C6073 XB2.XA1.MN0.D a_13808_1742# 1.71e-19
C6074 XB1.XA1.MN0.D XB1.XA3.MN0.S 0.00304f
C6075 XB1.XA4.MN0.D a_9560_2094# 0.0492f
C6076 SAR_IN a_12368_1742# 0.0505f
C6077 XB2.XA4.MN0.D XB2.XA4.MP0.D 0.00106f
C6078 XA3.XA4.MN0.D XA3.XA1.XA1.MN0.S 0.0145f
C6079 XA5.XA6.MP0.G a_12368_40932# 4.24e-19
C6080 XA20.XA3a.MN0.D XA4.XA1.XA4.MN1.D 0.0124f
C6081 XA1.XA1.XA5.MN2.D a_2288_44452# 0.158f
C6082 XA8.XA1.XA5.MN2.D a_19928_44804# 0.153f
C6083 XA1.XA6.MP0.G a_2288_40580# 5.5e-19
C6084 XA6.XA4.MN0.G a_16040_42692# 0.00224f
C6085 XA3.XA7.MP0.D a_8480_50788# 3.29e-19
C6086 a_12368_51492# a_12368_51140# 0.0109f
C6087 XA0.XA7.MP0.G a_n232_51140# 0.0661f
C6088 a_21080_53252# VREF 0.00386f
C6089 XA7.XA9.MN1.G a_18560_50436# 0.01f
C6090 AVDD a_n232_47620# 0.00125f
C6091 XA5.XA1.XA5.MN2.G XA6.XA1.XA5.MN2.G 1.58f
C6092 XA20.XA2a.MN0.D XA6.XA1.XA1.MP2.D 0.0102f
C6093 a_13520_43748# XA5.XA1.XA2.MP0.D 0.0686f
C6094 a_12368_43748# XA5.XA1.XA5.MP0.D 0.00176f
C6095 XA1.XA3.MN0.G XA1.XA1.XA1.MN0.D 0.00142f
C6096 EN a_22448_43396# 5.7e-20
C6097 D<0> VREF 1.29f
C6098 AVDD a_13520_44452# 0.00125f
C6099 D<5> a_7328_49380# 0.00891f
C6100 a_23600_50788# XA20.XA3.MN0.D 6.05e-20
C6101 D<1> XA3.XA4.MN0.D 0.0133f
C6102 D<2> XA6.XA4.MN0.D 0.203f
C6103 D<8> li_14804_29004# 3.5e-20
C6104 EN a_21080_40932# 0.00558f
C6105 a_17408_42692# XA7.XA1.XA4.MP0.D 0.00176f
C6106 XA2.XA6.MP0.G a_4808_46916# 7.76e-20
C6107 XA6.XA6.MP0.G a_14888_47268# 1.38e-19
C6108 D<7> a_4808_45860# 1.06e-19
C6109 XA6.XA1.XA5.MN2.G a_13520_45508# 2.31e-19
C6110 AVDD a_n232_41988# 0.00125f
C6111 XA0.XA4.MN0.D a_n232_47972# 0.0788f
C6112 VREF XA8.XA4.MN0.G 0.258f
C6113 XA4.XA4.MN0.D XA4.XA4.MN0.G 0.707f
C6114 a_3440_54308# XA2.XA11.MN1.G 6.78e-19
C6115 AVDD XA20.XA10.MN1.D 2.12f
C6116 XA6.XA1.XA1.MN0.S XA6.XA1.XA1.MN0.D 0.0743f
C6117 a_3440_41284# XA1.XA1.XA1.MN0.D 0.00224f
C6118 XA3.XA4.MN0.D a_8480_44804# 9.24e-20
C6119 VREF a_12368_44804# 0.0691f
C6120 XA4.XA6.MP0.G XA4.XA1.XA5.MN1.D 7.41e-19
C6121 XA4.XA1.XA5.MN2.G XA4.XA1.XA4.MN1.D 0.0131f
C6122 a_18560_47268# a_19928_47268# 8.89e-19
C6123 XA7.XA6.MP0.G EN 0.0712f
C6124 AVDD XB2.XA4.MN0.D 3.77e-19
C6125 XA3.XA4.MN0.G a_9848_46212# 2.2e-19
C6126 XA4.XA4.MN0.G a_8480_46212# 2.2e-19
C6127 XA20.XA9.MP0.D a_23600_52900# 0.0992f
C6128 XA4.XA10.MP0.D XA4.XA10.MP0.G 0.194f
C6129 CK_SAMPLE XA0.XA8.MP0.D 3.93e-19
C6130 AVDD XA5.XA1.XA5.MN2.G 5.46f
C6131 a_8408_3854# a_8408_3502# 0.0109f
C6132 XA2.XA6.MP0.G XA2.XA1.XA1.MN0.S 0.0143f
C6133 a_2288_45508# XA1.XA1.XA5.MN2.D 0.0675f
C6134 a_13520_45508# a_14888_45508# 8.89e-19
C6135 XA20.XA3a.MN0.D XA1.XA1.XA5.MP0.D 7.25e-19
C6136 XA6.XA6.MP0.G a_14888_41636# 7.76e-20
C6137 XA2.XA4.MN0.G a_4808_43396# 0.0104f
C6138 XA8.XA4.MN0.G XA8.XA1.XA5.MN0.D 0.0198f
C6139 XA0.XA6.MP2.G a_920_40580# 4.07e-20
C6140 XA4.XA1.XA5.MN2.G a_8480_40228# 1.34e-19
C6141 XA3.XA1.XA5.MN2.G a_9848_40228# 4.72e-19
C6142 D<4> a_11000_40932# 4.07e-20
C6143 SARN a_11000_1742# 0.0409f
C6144 XA7.XA3.MN0.G a_18560_44452# 0.0934f
C6145 AVDD a_23600_49028# 0.00154f
C6146 XA1.XA9.MN1.G D<7> 0.0378f
C6147 CK_SAMPLE a_8480_49380# 0.00139f
C6148 XA6.XA9.MN1.G a_16040_51140# 0.0222f
C6149 a_3440_51844# a_3440_51492# 0.0109f
C6150 XA5.XA7.MP0.D a_12368_51492# 0.0877f
C6151 XA20.XA10.MN1.D XA20.XA3.MN0.D 0.0573f
C6152 a_12368_52196# XA6.XA1.XA5.MN2.G 3.39e-19
C6153 li_9184_30648# li_9184_30036# 0.00271f
C6154 XDAC1.XC0.XRES8.B XDAC1.XC64b<1>.XRES8.B 6.7e-19
C6155 XA3.XA3.MN0.G a_9848_41988# 7.98e-19
C6156 SARN XDAC2.XC1.XRES4.B 13.9f
C6157 a_8480_44100# a_8480_43748# 0.0109f
C6158 a_19928_44100# XA8.XA1.XA5.MN1.D 0.00176f
C6159 EN XA6.XA1.XA5.MN1.D 0.0157f
C6160 XA6.XA1.XA5.MN2.D a_14888_43044# 5.1e-20
C6161 XA20.XA2a.MN0.D a_2288_42340# 0.00768f
C6162 XA0.XA6.MP2.G li_9184_23688# 3.5e-20
C6163 D<4> XA4.XA6.MN0.D 0.00148f
C6164 XA2.XA1.XA5.MN2.G a_2288_49732# 0.00457f
C6165 a_2288_51492# VREF 0.00396f
C6166 a_11000_50788# a_11000_50436# 0.0109f
C6167 a_22448_51140# XA20.XA3a.MN0.G 4.06e-20
C6168 AVDD a_13520_45508# 0.00131f
C6169 XDAC1.XC32a<0>.XRES4.B XDAC1.XC32a<0>.XRES8.B 0.471f
C6170 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES2.B 0.0136f
C6171 XA3.XA1.XA4.MP1.D XA3.XA1.XA4.MN1.D 0.00918f
C6172 XA0.XA4.MN0.D li_9184_12636# 1.76e-19
C6173 EN XA1.XA1.XA1.MN0.S 0.139f
C6174 XA8.XA1.XA5.MN2.G XA8.XA3.MN0.G 5.78e-19
C6175 D<7> a_3440_46916# 0.00249f
C6176 AVDD XA3.XA1.XA4.MP1.D 0.0913f
C6177 XA20.XA3.MN0.D a_23600_49028# 0.0765f
C6178 VREF a_21080_49380# 0.0167f
C6179 a_23600_49732# a_23600_49380# 0.0109f
C6180 XA0.XA6.MP0.G a_n232_47972# 6.28e-19
C6181 D<3> a_13520_47268# 3.18e-19
C6182 SARP XDAC1.XC64b<1>.XRES8.B 27.7f
C6183 a_18560_41636# a_19928_41636# 8.89e-19
C6184 XA2.XA6.MP0.G a_5960_44804# 5.5e-19
C6185 XA3.XA4.MN0.G a_8480_47268# 0.157f
C6186 XA2.XA1.XA5.MN2.G XA2.XA1.XA2.MP0.D 0.126f
C6187 VREF a_11000_45860# 0.0178f
C6188 XA3.XA4.MN0.D a_7328_45860# 9.15e-20
C6189 AVDD a_5960_40228# 0.467f
C6190 D<5> XA3.XA1.XA5.MN1.D 0.00185f
C6191 AVDD a_12368_52196# 0.37f
C6192 XA7.XA11.MN1.G a_17408_52900# 0.00273f
C6193 XA6.XA12.MP0.G a_16040_52900# 1.28e-19
C6194 a_3440_53252# a_4808_53252# 8.89e-19
C6195 CK_SAMPLE a_21080_52548# 0.00113f
C6196 XA3.XA11.MN1.G XA2.XA10.MP0.G 0.0024f
C6197 a_5960_40228# a_7328_40228# 8.89e-19
C6198 XA7.XA4.MN0.G a_17408_44100# 6.11e-19
C6199 XA1.XA4.MN0.G EN 0.0578f
C6200 XA0.XA4.MN0.G XA0.XA1.XA5.MN1.D 0.0242f
C6201 XA1.XA4.MN0.D a_3440_43044# 9.24e-20
C6202 XA6.XA1.XA5.MN2.G a_14888_41284# 0.0044f
C6203 XA0.XA11.MN1.G a_13808_n18# 0.00214f
C6204 a_7328_46212# a_7328_45860# 0.0109f
C6205 D<3> a_13520_41636# 6.49e-19
C6206 XA7.XA3.MN0.G a_18560_45508# 0.106f
C6207 XA1.XA3.MN0.G XA1.XA1.XA5.MN2.D 0.755f
C6208 XA20.XA10.MN1.D a_23600_50788# 0.0732f
C6209 a_11000_52900# XA5.XA1.XA5.MN2.G 1.06e-19
C6210 AVDD a_23600_50084# 0.00159f
C6211 a_920_52196# XA0.XA7.MP0.D 0.0658f
C6212 a_12368_52196# a_13520_52196# 0.00133f
C6213 CK_SAMPLE XA5.XA6.MN0.D 0.0676f
C6214 a_8408_686# a_8408_334# 0.0109f
C6215 a_9560_686# CK_SAMPLE_BSSW 0.0693f
C6216 a_12368_686# a_13808_686# 8e-19
C6217 XA20.XA2a.MN0.D a_9848_43044# 1.43e-19
C6218 XA3.XA4.MN0.G a_8480_41636# 6.69e-20
C6219 a_920_44452# a_920_44100# 0.0109f
C6220 a_3440_44804# EN 7.78e-19
C6221 XA7.XA6.MP0.G a_17408_39876# 0.00502f
C6222 XA1.XA4.MN0.D a_2288_40580# 9.15e-20
C6223 D<6> D<3> 0.0347f
C6224 a_21080_51140# D<0> 0.0672f
C6225 AVDD a_920_46564# 0.356f
C6226 a_8480_51140# a_8480_50788# 0.0109f
C6227 a_19928_51140# XA8.XA6.MN2.D 0.00176f
C6228 XA0.XA6.MP2.G D<1> 0.0959f
C6229 XA7.XA9.MN1.G a_17408_49732# 0.0215f
C6230 XA3.XA7.MP0.D a_8480_50084# 7.44e-20
C6231 D<5> D<4> 0.348f
C6232 D<7> D<2> 6.94e-19
C6233 XA2.XA1.XA5.MN2.G a_2288_50436# 0.0046f
C6234 XB2.XA3.MN1.D m3_16544_4532# 0.0137f
C6235 XA2.XA4.MN0.D li_9184_23688# 0.00504f
C6236 EN XA5.XA1.XA4.MP0.D 0.0386f
C6237 XA1.XA6.MP0.G XDAC2.XC32a<0>.XRES16.B 1.21e-19
C6238 XA5.XA6.MP0.G XDAC2.XC32a<0>.XRES4.B 0.00405f
C6239 XA20.XA2a.MN0.D a_8480_40580# 0.00123f
C6240 a_920_43396# a_920_43044# 0.0109f
C6241 a_23600_50084# XA20.XA3.MN0.D 0.00218f
C6242 a_11000_50084# a_11000_49732# 0.0109f
C6243 XA8.XA7.MP0.G a_21080_47972# 0.00363f
C6244 XA6.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.963f
C6245 D<3> a_12368_48324# 0.0164f
C6246 XA20.XA3.MN1.D a_23600_49732# 0.0137f
C6247 XA20.XA3a.MN0.G VREF 0.0339f
C6248 AVDD XA0.XA1.XA5.MP0.D 0.159f
C6249 SARP a_11000_1742# 0.00949f
C6250 D<8> XDAC2.XC128a<1>.XRES4.B 0.00406f
C6251 a_12368_42340# a_12368_41988# 0.0109f
C6252 a_n232_48324# a_n232_47972# 0.0109f
C6253 a_7328_48324# XA3.XA4.MN0.G 0.0674f
C6254 a_17408_48324# a_18560_48324# 0.00133f
C6255 XA5.XA1.XA5.MN2.G a_13520_44452# 5.11e-19
C6256 XA6.XA1.XA5.MN2.G a_12368_44452# 0.00486f
C6257 AVDD a_14888_41284# 0.00125f
C6258 XA2.XA6.MP0.G a_4808_45860# 7.76e-20
C6259 XA6.XA6.MP0.G a_14888_46212# 4.4e-19
C6260 AVDD a_9848_52900# 0.00166f
C6261 XA20.XA11.MN0.D XA20.XA9.MP0.D 0.0233f
C6262 DONE XA8.XA10.MP0.D 0.00436f
C6263 XA4.XA11.MN1.G a_11000_53604# 0.0658f
C6264 XA4.XA1.XA1.MN0.S a_9848_39876# 2.54e-19
C6265 XA4.XA1.XA1.MP1.D a_11000_40580# 0.00176f
C6266 a_n232_40932# a_n232_40580# 0.0109f
C6267 XA5.XA6.MP0.G a_12368_43396# 5.5e-19
C6268 a_920_46564# a_2288_46564# 8.89e-19
C6269 XA1.XA6.MP0.G a_2288_43044# 5.5e-19
C6270 XA4.XA4.MN0.G a_9848_45156# 0.00865f
C6271 XA4.XA3.MN0.G a_9848_46564# 0.156f
C6272 a_19928_46916# a_19928_46564# 0.0109f
C6273 XA8.XA7.MP0.G a_19928_42340# 3.12e-19
C6274 XA8.XA1.XA5.MN2.G a_21080_42340# 1.97e-19
C6275 XA2.XA1.XA5.MN2.G a_3440_41988# 0.0673f
C6276 XA0.XA4.MN0.D a_920_43748# 9.14e-20
C6277 XA6.XA10.MP0.G XA6.XA9.MN1.G 0.202f
C6278 AVDD a_22448_50788# 0.482f
C6279 CK_SAMPLE XA4.XA6.MN2.D 0.0389f
C6280 a_4808_52548# XA2.XA9.MN1.G 0.0727f
C6281 XB1.XA1.MP0.D XB1.XA3.MN0.S 6.58e-19
C6282 a_13808_2446# a_13808_2094# 0.0109f
C6283 XB1.M1.G a_11000_2094# 0.00148f
C6284 XB2.M1.G XB2.XA4.MP0.D 0.233f
C6285 D<2> a_16040_39876# 7.76e-20
C6286 SARN li_14804_29004# 0.00103f
C6287 XA20.XA3a.MN0.D XA3.XA1.XA4.MN1.D 0.0124f
C6288 a_8480_45156# a_8480_44804# 0.0109f
C6289 XA20.XA2a.MN0.D a_4808_43748# 4.48e-20
C6290 a_21080_45156# a_22448_45156# 8.89e-19
C6291 XA6.XA4.MN0.G a_14888_42692# 0.0049f
C6292 XA7.XA9.MN1.G a_17408_50436# 7.76e-19
C6293 AVDD XA20.XA3a.MN0.D 9.87f
C6294 XA20.XA10.MN1.D a_23600_49028# 0.00407f
C6295 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES2.B 0.0136f
C6296 XDAC2.X16ab.XRES4.B XDAC2.X16ab.XRES8.B 0.471f
C6297 XA20.XA2a.MN0.D XA6.XA1.XA1.MN0.S 0.137f
C6298 XA8.XA1.XA5.MP1.D XA8.XA1.XA5.MP0.D 0.0488f
C6299 XA4.XA1.XA5.MN1.D a_9848_43396# 0.00176f
C6300 EN a_21080_43396# 0.162f
C6301 a_23600_50436# XA20.XA3.MN1.D 0.00176f
C6302 AVDD a_12368_44452# 0.357f
C6303 XA2.XA1.XA5.MN2.G a_2288_48676# 0.00363f
C6304 D<1> XA2.XA4.MN0.D 3.88e-19
C6305 a_11000_50436# a_11000_50084# 0.0109f
C6306 XDAC2.XC64a<0>.XRES4.B XDAC2.XC1.XRES4.B 0.00284f
C6307 XDAC1.XC64a<0>.XRES16.B li_9184_9768# 0.00117f
C6308 XDAC2.XC64a<0>.XRES2.B XDAC2.XC64a<0>.XRES1A.B 0.0136f
C6309 li_14804_10380# li_14804_9768# 0.00271f
C6310 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES4.B 0.00405f
C6311 XA3.XA1.XA2.MP0.D a_7328_41284# 1.07e-19
C6312 XA6.XA1.XA4.MP1.D a_16040_42340# 0.00176f
C6313 a_4808_42692# a_4808_42340# 0.0109f
C6314 D<3> a_13520_46212# 0.0141f
C6315 a_11000_49028# a_11000_48676# 0.0109f
C6316 XA20.XA3.MN0.D XA20.XA3a.MN0.D 0.176f
C6317 D<7> a_3440_45860# 0.0675f
C6318 XA6.XA1.XA5.MN2.G a_12368_45508# 0.00595f
C6319 XA5.XA1.XA5.MN2.G a_13520_45508# 9.01e-20
C6320 AVDD a_23600_42340# 0.00405f
C6321 VREF XA7.XA4.MN0.G 0.263f
C6322 XA3.XA4.MN0.D XA4.XA4.MN0.G 3.16e-20
C6323 XA4.XA4.MN0.D XA3.XA4.MN0.G 3.16e-20
C6324 a_2288_54308# XA2.XA11.MN1.G 8.3e-19
C6325 AVDD XA8.XA12.MP0.G 0.71f
C6326 a_14888_54308# a_14888_53956# 0.0109f
C6327 a_920_53956# a_2288_53956# 8.89e-19
C6328 SARP li_9184_18564# 0.00103f
C6329 XA1.XA1.XA1.MP2.D a_2288_40932# 0.00176f
C6330 a_14888_41284# a_16040_41284# 0.00133f
C6331 XA3.XA4.MN0.D a_7328_44804# 9.15e-20
C6332 VREF a_11000_44804# 0.0691f
C6333 D<4> a_11000_43396# 7.76e-20
C6334 XA4.XA1.XA5.MN2.G XA3.XA1.XA4.MN1.D 7.2e-19
C6335 XA0.XA6.MP2.G a_920_43044# 7.76e-20
C6336 a_5960_47268# a_5960_46916# 0.0109f
C6337 XA0.XA6.MP0.G a_920_43748# 5.5e-19
C6338 AVDD XB2.M1.G 0.717f
C6339 XA3.XA4.MN0.G a_8480_46212# 0.0149f
C6340 XA20.XA9.MP0.D a_22448_52900# 0.0026f
C6341 a_9848_52900# a_11000_52900# 0.00133f
C6342 CK_SAMPLE a_23600_51844# 7.93e-19
C6343 AVDD XA4.XA1.XA5.MN2.G 4.81f
C6344 XA3.XA11.MN1.G XA3.XA7.MP0.D 0.00283f
C6345 XA7.XA11.MN1.G a_18560_52196# 5.56e-19
C6346 a_8408_3854# a_9560_3854# 0.00133f
C6347 XA20.XA3a.MN0.D XA1.XA1.XA2.MP0.D 0.199f
C6348 XA8.XA4.MN0.G XA8.XA1.XA2.MP0.D 0.206f
C6349 XA0.XA6.MP2.G a_n232_40580# 5.24e-19
C6350 XA3.XA1.XA5.MN2.G a_8480_40228# 0.0825f
C6351 XA4.XA1.XA5.MN2.G a_7328_40228# 0.00255f
C6352 D<4> a_9848_40932# 5.24e-19
C6353 SARN a_9560_1742# 2.97e-20
C6354 XA20.XA3.MN0.D a_23600_42340# 2.14e-19
C6355 D<8> a_920_44100# 0.00245f
C6356 XA7.XA3.MN0.G a_17408_44452# 0.055f
C6357 AVDD a_22448_49028# 0.488f
C6358 CK_SAMPLE a_7328_49380# 7.89e-19
C6359 XA6.XA9.MN1.G a_14888_51140# 0.0469f
C6360 a_11000_51844# XA4.XA8.MP0.D 0.0215f
C6361 a_19928_51844# a_21080_51844# 0.00133f
C6362 XA20.XA10.MN1.D a_23600_50084# 0.0046f
C6363 a_17408_53956# VREF 0.00396f
C6364 D<5> XDAC1.X16ab.XRES8.B 1.85e-19
C6365 EN XA5.XA1.XA5.MN1.D 0.0157f
C6366 XA20.XA2a.MN0.D a_920_42340# 0.00732f
C6367 XA3.XA3.MN0.G a_8480_41988# 0.00343f
C6368 D<4> XA4.XA6.MP0.G 2.1f
C6369 XA0.XA7.MP0.G a_2288_49732# 7.1e-20
C6370 XA2.XA1.XA5.MN2.G a_920_49732# 7.1e-20
C6371 a_920_51492# VREF 0.00396f
C6372 D<3> XA3.XA6.MP0.G 0.0672f
C6373 D<1> XA1.XA6.MP0.G 0.037f
C6374 D<2> XA2.XA6.MP0.G 0.0297f
C6375 AVDD a_12368_45508# 0.359f
C6376 a_22448_50788# a_23600_50788# 0.00133f
C6377 XA8.XA1.XA2.MP0.D XA8.XA1.XA4.MP0.D 4.34e-19
C6378 a_19928_43044# XA8.XA1.XA4.MN1.D 0.00176f
C6379 a_8480_43044# a_8480_42692# 0.0109f
C6380 XA8.XA1.XA5.MN2.G XA7.XA3.MN0.G 0.106f
C6381 D<7> a_2288_46916# 0.0185f
C6382 AVDD XA2.XA1.XA4.MP1.D 0.0913f
C6383 a_3440_49380# a_4808_49380# 8.89e-19
C6384 XA5.XA4.MN0.D a_13520_49380# 0.155f
C6385 VREF a_19928_49380# 8.08e-19
C6386 XA2.XA6.MP0.G XA2.XA4.MN0.G 0.0408f
C6387 XA20.XA3.MN1.D a_23600_48676# 0.0604f
C6388 D<3> a_12368_47268# 0.0148f
C6389 a_5960_41636# XA2.XA1.XA1.MP2.D 0.00176f
C6390 XA2.XA6.MP0.G a_4808_44804# 7.76e-20
C6391 D<1> a_18560_44100# 6.49e-19
C6392 a_12368_47972# a_12368_47620# 0.0109f
C6393 XA6.XA6.MP0.G a_16040_45156# 5.5e-19
C6394 XA3.XA4.MN0.G a_7328_47268# 0.155f
C6395 XA8.XA7.MP0.G a_22448_43748# 0.00113f
C6396 XA0.XA7.MP0.G XA2.XA1.XA2.MP0.D 1.74e-19
C6397 XA2.XA1.XA5.MN2.G XA1.XA1.XA5.MN0.D 7.2e-19
C6398 VREF a_9848_45860# 1.19e-19
C6399 AVDD a_4808_40228# 0.00131f
C6400 D<5> XA3.XA1.XA5.MP1.D 7.43e-19
C6401 AVDD a_11000_52196# 0.37f
C6402 XA7.XA11.MN1.G a_16040_52900# 0.00183f
C6403 XA6.XA12.MP0.G a_14888_52900# 0.00258f
C6404 DONE SARN 3.94e-19
C6405 XA5.XA11.MP0.D a_12368_53252# 0.0494f
C6406 CK_SAMPLE a_19928_52548# 3.41e-19
C6407 a_13520_53604# XA5.XA10.MP0.D 1.17e-19
C6408 a_22448_53604# a_22448_53252# 0.0109f
C6409 a_18560_40580# a_18560_40228# 0.0109f
C6410 D<7> XA1.XA1.XA1.MN0.S 0.0133f
C6411 XA0.XA4.MN0.G EN 0.227f
C6412 XA1.XA4.MN0.D a_2288_43044# 9.15e-20
C6413 XA6.XA1.XA5.MN2.G a_13520_41284# 0.00733f
C6414 XA0.XA11.MN1.G a_12368_n18# 0.00164f
C6415 XA20.XA3a.MN0.D a_13520_44452# 2.59e-20
C6416 a_18560_46212# a_19928_46212# 8.89e-19
C6417 D<3> a_12368_41636# 7.77e-20
C6418 XA7.XA3.MN0.G a_17408_45508# 0.0682f
C6419 XA6.XA9.MN0.D XA6.XA7.MP0.D 0.00986f
C6420 XA4.XA10.MP0.G a_9848_51492# 6.8e-20
C6421 XA20.XA10.MN1.D a_22448_50788# 0.0674f
C6422 AVDD a_22448_50084# 0.366f
C6423 a_n232_52196# XA0.XA7.MP0.D 0.0678f
C6424 CK_SAMPLE XA5.XA6.MP0.D 0.0278f
C6425 a_8408_686# CK_SAMPLE_BSSW 0.0674f
C6426 a_12368_44452# a_13520_44452# 0.00133f
C6427 XA20.XA2a.MN0.D a_8480_43044# 1.43e-19
C6428 XA4.XA1.XA5.MN2.D a_11000_43748# 0.00388f
C6429 XA20.XA3a.MN0.D a_n232_41988# 0.00542f
C6430 a_2288_44804# EN 3.4e-19
C6431 XA7.XA6.MP0.G a_16040_39876# 0.00308f
C6432 SARN XDAC2.XC128a<1>.XRES4.B 13.9f
C6433 D<5> XA3.XA6.MN2.D 1.59e-19
C6434 AVDD a_n232_46564# 0.00125f
C6435 XA8.XA1.XA5.MN2.G a_18560_50788# 1.87e-19
C6436 XA2.XA1.XA5.MN2.G a_920_50436# 7.1e-20
C6437 XA0.XA7.MP0.G a_2288_50436# 7.1e-20
C6438 XA2.XA9.MN1.G XA2.XA4.MN0.D 0.00938f
C6439 XA3.XA9.MN1.G VREF 0.0732f
C6440 XA20.XA10.MN1.D XA20.XA3a.MN0.D 0.0141f
C6441 XB2.XA3.MN1.D m3_16472_4532# 0.0137f
C6442 XDAC1.XC128b<2>.XRES16.B XDAC1.XC128b<2>.XRES1A.B 0.454f
C6443 XDAC2.XC128b<2>.XRES16.B li_14804_20208# 0.00117f
C6444 XA3.XA4.MN0.D XDAC1.X16ab.XRES16.B 0.00136f
C6445 XA0.XA6.MP0.G li_14804_13248# 1.85e-20
C6446 EN XA4.XA1.XA4.MP0.D 0.0386f
C6447 XA5.XA1.XA5.MN0.D a_13520_43044# 0.00176f
C6448 a_12368_43396# a_13520_43396# 0.00133f
C6449 XA5.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.885f
C6450 XA20.XA3.MN6.D a_23600_49732# 8.29e-20
C6451 XA20.XA3.MN1.D a_22448_49732# 8.29e-20
C6452 XA8.XA6.MP0.D VREF 0.0146f
C6453 D<7> XA1.XA4.MN0.G 0.259f
C6454 AVDD XA0.XA1.XA5.MN0.D 0.00889f
C6455 XA2.XA1.XA5.MN2.G a_2288_47620# 0.00363f
C6456 SARP a_9560_1742# 9.76e-19
C6457 XA6.XA1.XA5.MN2.G a_11000_44452# 7.1e-20
C6458 XA5.XA1.XA5.MN2.G a_12368_44452# 7.1e-20
C6459 D<7> a_3440_44804# 5.26e-19
C6460 XA20.XA10.MN1.D a_23600_42340# 0.00431f
C6461 AVDD a_13520_41284# 0.00125f
C6462 XA2.XA4.MN0.D a_5960_46916# 0.00254f
C6463 AVDD a_8480_52900# 0.00166f
C6464 a_21080_53956# a_21080_53604# 0.0109f
C6465 XA3.XA12.MP0.G a_8480_53604# 0.102f
C6466 XA4.XA11.MN1.G a_9848_53604# 0.0709f
C6467 SARP XDAC1.XC1.XRES4.B 13.9f
C6468 XA4.XA1.XA1.MN0.D a_11000_40580# 8.3e-19
C6469 a_11000_40932# a_12368_40932# 8.89e-19
C6470 XA3.XA4.MN0.G a_9848_45156# 2.2e-19
C6471 XA4.XA4.MN0.G a_8480_45156# 2.2e-19
C6472 XA8.XA1.XA5.MN2.G a_19928_42340# 0.00568f
C6473 XA0.XA7.MP0.G a_3440_41988# 0.0039f
C6474 XA2.XA1.XA5.MN2.G a_2288_41988# 0.0734f
C6475 XA0.XA4.MN0.D a_n232_43748# 9.25e-20
C6476 VREF XA8.XA1.XA5.MP1.D 0.00623f
C6477 a_16040_52548# a_17408_52548# 8.89e-19
C6478 XA20.XA9.MP0.D a_23600_52196# 0.0037f
C6479 AVDD a_21080_50788# 0.361f
C6480 CK_SAMPLE D<4> 0.0523f
C6481 XB2.M1.G XB2.XA4.MN0.D 0.139f
C6482 XB1.M1.G a_9560_2094# 0.0193f
C6483 XB1.XA4.MP0.D a_8408_2094# 0.0682f
C6484 D<2> a_14888_39876# 0.00212f
C6485 XA20.XA3a.MN0.D XA3.XA1.XA4.MP1.D 0.0124f
C6486 XA0.XA1.XA5.MN2.D a_920_44452# 0.158f
C6487 XA7.XA1.XA5.MN2.D a_18560_44804# 0.153f
C6488 XA20.XA2a.MN0.D a_3440_43748# 2.91e-20
C6489 XA3.XA3.MN0.G XA3.XA1.XA2.MP0.D 0.0363f
C6490 a_11000_51492# a_11000_51140# 0.0109f
C6491 XA20.XA4.MN0.D XA20.XA3.MN6.D 0.0887f
C6492 AVDD a_23600_47972# 0.00159f
C6493 XA1.XA9.MN1.G XA1.XA6.MN0.D 0.0615f
C6494 XA20.XA10.MN1.D a_22448_49028# 1.78e-19
C6495 XA4.XA1.XA5.MN2.G XA5.XA1.XA5.MN2.G 0.0255f
C6496 XA20.XA2a.MN0.D XA5.XA1.XA1.MP2.D 0.0102f
C6497 XA3.XA6.MP0.G li_14804_24912# 0.00504f
C6498 XA1.XA6.MP0.G XDAC2.X16ab.XRES16.B 1.21e-19
C6499 EN a_19928_43396# 0.00238f
C6500 XA3.XA6.MP0.G XA6.XA6.MP0.G 0.0273f
C6501 XA2.XA6.MP0.G XA7.XA6.MP0.G 0.0311f
C6502 XA4.XA6.MP0.G XA5.XA6.MP0.G 6.62f
C6503 a_23600_50436# XA20.XA3.MN6.D 0.0215f
C6504 AVDD a_11000_44452# 0.357f
C6505 XA0.XA7.MP0.G a_2288_48676# 7.1e-20
C6506 XA2.XA1.XA5.MN2.G a_920_48676# 7.1e-20
C6507 D<1> XA1.XA4.MN0.D 0.0342f
C6508 XA7.XA6.MP2.D VREF 5.13e-19
C6509 D<8> XDAC2.XC64b<1>.XRES4.B 4.06e-21
C6510 a_16040_42692# XA6.XA1.XA4.MP0.D 0.00176f
C6511 D<3> a_12368_46212# 0.0202f
C6512 a_22448_49028# a_23600_49028# 0.00133f
C6513 XA20.XA3.MN0.D a_23600_47972# 0.0329f
C6514 D<7> a_2288_45860# 0.0774f
C6515 XA5.XA1.XA5.MN2.G a_12368_45508# 7.1e-20
C6516 XA6.XA1.XA5.MN2.G a_11000_45508# 7.1e-20
C6517 AVDD a_22448_42340# 0.575f
C6518 VREF XA6.XA4.MN0.G 0.263f
C6519 XA3.XA4.MN0.D XA3.XA4.MN0.G 0.728f
C6520 a_3440_54308# XA0.XA12.MP0.D 0.00123f
C6521 AVDD XA7.XA12.MP0.G 0.706f
C6522 a_2288_41284# XA1.XA1.XA1.MP1.D 0.00176f
C6523 XA1.XA1.XA1.MN0.S a_2288_40932# 0.0271f
C6524 XA4.XA1.XA5.MN2.G XA3.XA1.XA4.MP1.D 0.00353f
C6525 XA3.XA1.XA5.MN2.G XA3.XA1.XA4.MN1.D 0.0131f
C6526 XA0.XA6.MP2.G a_n232_43044# 6.49e-19
C6527 a_17408_47268# a_18560_47268# 0.00133f
C6528 AVDD XB1.XA4.MN0.D 3.77e-19
C6529 VREF a_9848_44804# 7.12e-19
C6530 D<4> a_9848_43396# 6.49e-19
C6531 XA0.XA6.MP0.G a_n232_43748# 7.76e-20
C6532 XA3.XA4.MN0.G a_7328_46212# 3.46e-19
C6533 XA3.XA10.MP0.D XA3.XA10.MP0.G 0.194f
C6534 CK_SAMPLE a_22448_51844# 0.00684f
C6535 AVDD XA3.XA1.XA5.MN2.G 5.46f
C6536 XA3.XA11.MN1.G XA2.XA7.MP0.D 8.25e-19
C6537 XA7.XA11.MN1.G a_17408_52196# 7.34e-19
C6538 a_920_45508# XA0.XA1.XA5.MN2.D 0.0659f
C6539 a_12368_45508# a_13520_45508# 0.00133f
C6540 a_17408_45860# XA7.XA1.XA5.MN2.D 3.12e-20
C6541 XA20.XA3a.MN0.D XA0.XA1.XA5.MP0.D 7.08e-19
C6542 XA1.XA4.MN0.G a_3440_43396# 0.0104f
C6543 XA3.XA1.XA5.MN2.G a_7328_40228# 0.0128f
C6544 D<8> a_n232_44100# 0.00767f
C6545 AVDD a_21080_49028# 0.356f
C6546 CK_SAMPLE a_5960_49380# 7.89e-19
C6547 XA6.XA9.MN1.G a_13520_51140# 2.84e-19
C6548 a_2288_51844# a_2288_51492# 0.0109f
C6549 a_9848_51844# XA4.XA8.MP0.D 0.0215f
C6550 XA4.XA7.MP0.D a_11000_51492# 0.0893f
C6551 a_16040_53956# VREF 0.00366f
C6552 a_11000_52196# XA5.XA1.XA5.MN2.G 3.39e-19
C6553 XDAC2.XC0.XRES16.B XDAC2.XC0.XRES1A.B 0.454f
C6554 a_7328_44100# a_7328_43748# 0.0109f
C6555 a_18560_44100# XA7.XA1.XA5.MN1.D 0.00176f
C6556 EN XA5.XA1.XA5.MP1.D 0.0543f
C6557 XA2.XA1.XA5.MN1.D XA2.XA1.XA5.MP1.D 0.00918f
C6558 XA20.XA3a.MN0.D a_14888_41284# 0.00649f
C6559 XA5.XA1.XA5.MN2.D a_13520_43044# 5.1e-20
C6560 XA20.XA2a.MN0.D a_n232_42340# 0.0843f
C6561 XA0.XA6.MP2.G XDAC1.X16ab.XRES16.B 3.84e-19
C6562 SARN li_14804_8736# 0.00103f
C6563 XA8.XA6.MP2.D a_21080_50436# 0.00176f
C6564 a_9848_50788# a_9848_50436# 0.0109f
C6565 XA0.XA7.MP0.G a_920_49732# 0.00457f
C6566 AVDD a_11000_45508# 0.359f
C6567 li_14804_15696# li_14804_15084# 0.00271f
C6568 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES8.B 0.0228f
C6569 XDAC2.XC128a<1>.XRES16.B XDAC2.XC32a<0>.XRES16.B 0.0114f
C6570 XA0.XA1.XA2.MP0.D a_920_41988# 0.0219f
C6571 XA4.XA1.XA2.MP0.D a_11000_42340# 2.54e-19
C6572 XA8.XA1.XA2.MP0.D XA8.XA1.XA4.MN0.D 0.056f
C6573 XA1.XA4.MN0.D XDAC1.XC32a<0>.XRES16.B 1.21e-19
C6574 XA0.XA4.MN0.D li_9184_13248# 1.85e-20
C6575 EN XA0.XA1.XA1.MN0.S 0.17f
C6576 AVDD XA2.XA1.XA4.MN1.D 0.00889f
C6577 XA8.XA1.XA5.MN2.G XA6.XA3.MN0.G 6.95e-19
C6578 XA7.XA1.XA5.MN2.G XA7.XA3.MN0.G 0.00127f
C6579 XA5.XA4.MN0.D a_12368_49380# 0.154f
C6580 a_22448_49732# a_22448_49380# 0.0109f
C6581 VREF a_18560_49380# 8.08e-19
C6582 XA20.XA9.MP0.D a_23600_44452# 0.00334f
C6583 XA20.XA3.MN1.D a_22448_48676# 0.0526f
C6584 XA20.XA3.MN6.D a_23600_48676# 5.18e-19
C6585 a_17408_41636# a_18560_41636# 0.00133f
C6586 a_5960_41636# XA2.XA1.XA1.MN0.S 0.0694f
C6587 SARP li_9184_29004# 0.00103f
C6588 XA6.XA6.MP0.G a_14888_45156# 7.76e-20
C6589 XA8.XA7.MP0.G a_21080_43748# 0.00442f
C6590 D<3> EN 0.0683f
C6591 XA2.XA1.XA5.MN2.G XA1.XA1.XA5.MP0.D 0.00353f
C6592 XA2.XA4.MN0.D a_5960_45860# 9.14e-20
C6593 VREF a_8480_45860# 1.19e-19
C6594 AVDD a_3440_40228# 0.00131f
C6595 D<1> a_17408_44100# 7.77e-20
C6596 XA2.XA11.MN1.G XA2.XA10.MP0.G 7.66e-19
C6597 AVDD a_9848_52196# 0.00154f
C6598 DONE XA8.XA9.MN0.D 0.00105f
C6599 a_2288_53252# a_3440_53252# 0.00133f
C6600 a_4808_40228# a_5960_40228# 0.00133f
C6601 XA6.XA1.XA5.MN2.G a_12368_41284# 0.0169f
C6602 XA5.XA1.XA5.MN2.G a_13520_41284# 0.00392f
C6603 XA6.XA4.MN0.G a_16040_44100# 6.11e-19
C6604 XA7.XA6.MP0.G a_18560_42692# 7.76e-20
C6605 XA0.XA11.MN1.G a_11000_n18# 0.00164f
C6606 a_5960_46212# a_5960_45860# 0.0109f
C6607 XA3.XA6.MP0.G XA3.XA1.XA4.MN0.D 6.07e-19
C6608 D<8> XA0.XA1.XA5.MN2.D 0.753f
C6609 XA6.XA9.MN1.G XA6.XA7.MP0.D 0.274f
C6610 AVDD a_21080_50084# 0.361f
C6611 XA2.XA9.MN0.D a_4808_51844# 0.00176f
C6612 XA2.XA9.MN1.G a_5960_51844# 6.57e-19
C6613 CK_SAMPLE XA5.XA6.MP0.G 0.0463f
C6614 a_11000_52196# a_12368_52196# 8.89e-19
C6615 a_11000_686# a_12368_686# 8.89e-19
C6616 XB2.XA3.MN1.D a_14960_n18# 0.0124f
C6617 XA4.XA1.XA5.MN2.D a_9848_43748# 0.00224f
C6618 a_n232_44452# a_n232_44100# 0.0109f
C6619 a_920_44804# EN 3.4e-19
C6620 XA7.XA6.MP0.G a_14888_39876# 0.00296f
C6621 D<5> XA3.XA6.MP2.D 0.0399f
C6622 a_7328_51140# a_7328_50788# 0.0109f
C6623 XA8.XA1.XA5.MN2.G a_17408_50788# 0.00548f
C6624 AVDD XA8.XA3.MN0.G 2.49f
C6625 a_920_51492# XA0.XA6.MP0.G 4.06e-20
C6626 XA0.XA7.MP0.G a_920_50436# 0.0046f
C6627 XA20.XA10.MN1.D a_23600_47972# 0.00517f
C6628 XB2.XA4.MP0.D m3_16544_308# 0.0634f
C6629 EN XA4.XA1.XA4.MN0.D 3.17e-19
C6630 a_n232_43396# a_n232_43044# 0.0109f
C6631 XA2.XA4.MN0.D XDAC1.X16ab.XRES16.B 0.0181f
C6632 a_22448_50084# a_23600_50084# 0.00133f
C6633 a_9848_50084# a_9848_49732# 0.0109f
C6634 XA4.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.963f
C6635 XA3.XA6.MP0.G a_8480_49380# 0.0547f
C6636 XA20.XA3.MN6.D a_22448_49732# 0.0157f
C6637 XA20.XA9.MP0.D a_23600_45508# 0.00334f
C6638 AVDD XA0.XA1.XA2.MP0.D 0.263f
C6639 XA0.XA7.MP0.G a_2288_47620# 7.1e-20
C6640 XA2.XA1.XA5.MN2.G a_920_47620# 7.1e-20
C6641 a_11000_42340# a_11000_41988# 0.0109f
C6642 XA20.XA1.MN0.D a_23600_41988# 0.056f
C6643 a_11000_42692# XA4.XA1.XA1.MN0.S 6.76e-20
C6644 D<8> li_14804_19176# 0.00508f
C6645 XA5.XA1.XA5.MN2.G a_11000_44452# 0.00486f
C6646 D<7> a_2288_44804# 2.37e-19
C6647 a_5960_48324# XA2.XA4.MN0.G 0.0658f
C6648 a_16040_48324# a_17408_48324# 8.89e-19
C6649 AVDD a_12368_41284# 0.361f
C6650 VREF a_7328_46916# 0.0536f
C6651 XA2.XA4.MN0.D a_4808_46916# 0.00456f
C6652 D<3> a_13520_45156# 7.77e-19
C6653 AVDD a_7328_52900# 0.387f
C6654 XA3.XA12.MP0.G a_7328_53604# 0.0877f
C6655 XA4.XA11.MN1.G a_8480_53604# 0.00787f
C6656 XA4.XA1.XA1.MN0.D a_9848_40580# 0.035f
C6657 XA0.XA11.MN1.G a_13808_3150# 0.0101f
C6658 a_n232_46564# a_920_46564# 0.00133f
C6659 XA3.XA4.MN0.G a_8480_45156# 0.00865f
C6660 XA3.XA3.MN0.G a_8480_46564# 0.156f
C6661 a_18560_46916# a_18560_46564# 0.0109f
C6662 XA8.XA1.XA5.MN2.G a_18560_42340# 4.69e-19
C6663 XA5.XA10.MP0.G XA5.XA9.MN0.D 0.106f
C6664 a_3440_52548# XA1.XA9.MN0.D 0.00176f
C6665 AVDD a_19928_50788# 0.00154f
C6666 CK_SAMPLE XA3.XA6.MN2.D 0.0389f
C6667 a_12368_2446# a_12368_2094# 0.0109f
C6668 SAR_IP a_11000_1742# 0.0505f
C6669 XB1.M1.G a_8408_2094# 0.0982f
C6670 XB2.XA1.MP0.D XB2.XA0.MP0.D 0.0524f
C6671 XA2.XA4.MN0.D XA2.XA1.XA1.MN0.S 0.0163f
C6672 D<2> a_13520_39876# 1.27e-19
C6673 SARN XDAC2.XC64b<1>.XRES4.B 13.9f
C6674 XA20.XA3a.MN0.D XA2.XA1.XA4.MP1.D 0.0124f
C6675 XA0.XA1.XA5.MN2.D a_n232_44452# 0.153f
C6676 XA7.XA1.XA5.MN2.D a_17408_44804# 0.156f
C6677 a_7328_45156# a_7328_44804# 0.0109f
C6678 a_19928_45156# a_21080_45156# 0.00133f
C6679 XA5.XA4.MN0.G a_13520_42692# 0.0049f
C6680 a_17408_53252# VREF 0.00267f
C6681 XA20.XA4.MN0.D XA20.XA3a.MN0.G 0.00384f
C6682 AVDD a_22448_47972# 0.389f
C6683 a_12368_51844# D<3> 1.25e-19
C6684 XA1.XA9.MN1.G XA1.XA6.MP0.D 0.0618f
C6685 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES2.B 0.0136f
C6686 XDAC1.X16ab.XRES4.B XDAC1.X16ab.XRES8.B 0.471f
C6687 a_11000_43748# XA4.XA1.XA5.MP0.D 0.00176f
C6688 XA3.XA1.XA5.MN1.D a_8480_43396# 0.00176f
C6689 XA0.XA1.XA5.MN0.D XA0.XA1.XA5.MP0.D 0.00918f
C6690 XA8.XA1.XA5.MN1.D XA8.XA1.XA5.MN0.D 0.0488f
C6691 XA8.XA1.XA5.MP1.D XA8.XA1.XA2.MP0.D 6.52e-20
C6692 XA20.XA2a.MN0.D XA5.XA1.XA1.MN0.S 0.137f
C6693 EN a_18560_43396# 0.00238f
C6694 XA0.XA7.MP0.G a_920_48676# 0.00363f
C6695 AVDD a_9848_44452# 0.00125f
C6696 a_23600_50436# XA20.XA3a.MN0.G 0.0658f
C6697 a_22448_50436# XA20.XA3.MN6.D 0.00322f
C6698 XA8.XA1.XA5.MN2.G a_17408_49028# 0.00363f
C6699 D<1> VREF 1.3f
C6700 D<2> XA3.XA4.MN0.D 0.0185f
C6701 a_9848_50436# a_9848_50084# 0.0109f
C6702 XA4.XA6.MP0.G XA4.XA6.MP0.D 0.0392f
C6703 XDAC1.XC64a<0>.XRES4.B XDAC1.XC1.XRES4.B 0.00284f
C6704 li_9184_10380# li_9184_9768# 0.00271f
C6705 XDAC1.XC64a<0>.XRES2.B XDAC1.XC64a<0>.XRES1A.B 0.0136f
C6706 XA1.XA3.MN0.G li_14804_29616# 0.00504f
C6707 EN a_17408_40932# 0.00564f
C6708 XA1.XA1.XA4.MP0.D XA1.XA1.XA4.MN0.D 0.00918f
C6709 XA6.XA1.XA4.MN1.D a_14888_42340# 0.00176f
C6710 a_3440_42692# a_3440_42340# 0.0109f
C6711 XA20.XA3.MN6.D a_23600_47620# 5.92e-19
C6712 a_9848_49028# a_9848_48676# 0.0109f
C6713 XA20.XA3.MN0.D a_22448_47972# 0.0218f
C6714 XA5.XA1.XA5.MN2.G a_11000_45508# 0.00595f
C6715 AVDD a_21080_42340# 0.361f
C6716 VREF XA5.XA4.MN0.G 0.263f
C6717 XA8.XA4.MN0.D a_21080_48324# 0.0698f
C6718 a_2288_54308# XA0.XA12.MP0.D 8.45e-19
C6719 AVDD XA8.XA11.MN1.G 1.04f
C6720 a_13520_54308# a_13520_53956# 0.0109f
C6721 a_n232_53956# a_920_53956# 0.00133f
C6722 SARP XDAC1.XC128a<1>.XRES4.B 13.9f
C6723 a_13520_41284# a_14888_41284# 8.89e-19
C6724 XA5.XA1.XA1.MN0.S XA5.XA1.XA1.MN0.D 0.0743f
C6725 XA5.XA1.XA1.MP2.D XA5.XA1.XA1.MP1.D 0.0488f
C6726 XA3.XA1.XA5.MN2.G XA3.XA1.XA4.MP1.D 7.44e-19
C6727 a_4808_47268# a_4808_46916# 0.0109f
C6728 VREF a_8480_44804# 7.12e-19
C6729 XA2.XA4.MN0.D a_5960_44804# 9.14e-20
C6730 XA6.XA6.MP0.G EN 0.0711f
C6731 AVDD XB1.XA4.MP0.D 2.39f
C6732 a_8480_52900# a_9848_52900# 8.89e-19
C6733 XA8.XA10.MP0.D a_21080_52900# 0.0893f
C6734 CK_SAMPLE a_21080_51844# 0.00182f
C6735 AVDD XA2.XA1.XA5.MN2.G 4.81f
C6736 XA7.XA11.MN1.G a_16040_52196# 4.29e-19
C6737 XA20.XA3a.MN0.D XA0.XA1.XA5.MN0.D 0.0106f
C6738 SARN XB2.XA0.MP0.D 0.00703f
C6739 a_n232_45508# XA0.XA1.XA5.MN2.D 0.0674f
C6740 XA1.XA4.MN0.G a_2288_43396# 8.07e-19
C6741 XA7.XA4.MN0.G XA7.XA1.XA5.MN0.D 0.0198f
C6742 XA3.XA1.XA5.MN2.G a_5960_40228# 0.0108f
C6743 D<1> XA7.XA1.XA1.MN0.D 0.0166f
C6744 XA6.XA3.MN0.G a_16040_44452# 0.055f
C6745 XA5.XA9.MN1.G a_14888_51140# 2.84e-19
C6746 AVDD a_19928_49028# 0.00154f
C6747 XA0.XA9.MN1.G XA0.XA6.MP2.D 0.0618f
C6748 CK_SAMPLE a_4808_49380# 0.00139f
C6749 a_18560_51844# a_19928_51844# 8.89e-19
C6750 XA4.XA7.MP0.D a_9848_51492# 0.124f
C6751 D<5> li_9184_25524# 0.00504f
C6752 EN XA4.XA1.XA5.MP1.D 0.0544f
C6753 XA20.XA3a.MN0.D a_13520_41284# 0.00649f
C6754 XA20.XA2a.MN0.D XA20.XA1.MN0.D 0.0119f
C6755 XA5.XA1.XA5.MN2.D a_12368_43044# 1.88e-19
C6756 XA8.XA1.XA5.MN2.G a_17408_50084# 0.00366f
C6757 XA7.XA8.MP0.D VREF 7.83e-19
C6758 AVDD a_9848_45508# 0.00131f
C6759 a_21080_50788# a_22448_50788# 8.89e-19
C6760 a_7328_43044# a_7328_42692# 0.0109f
C6761 a_18560_43044# XA7.XA1.XA4.MN1.D 0.00176f
C6762 XA4.XA1.XA2.MP0.D a_9848_42340# 0.095f
C6763 XA0.XA1.XA2.MP0.D a_n232_41988# 0.0568f
C6764 AVDD XA1.XA1.XA4.MN1.D 0.00889f
C6765 XA7.XA1.XA5.MN2.G XA6.XA3.MN0.G 0.106f
C6766 XA2.XA1.XA5.MN2.G a_2288_46564# 0.00363f
C6767 VREF a_17408_49380# 0.0171f
C6768 XA5.XA6.MP0.G a_13520_48324# 0.00295f
C6769 XA20.XA3.MN6.D a_22448_48676# 0.00982f
C6770 a_2288_49380# a_3440_49380# 0.00133f
C6771 a_17408_41988# XA7.XA1.XA1.MN0.S 3.8e-19
C6772 a_4808_41636# XA2.XA1.XA1.MN0.S 0.0674f
C6773 a_11000_47972# a_11000_47620# 0.0109f
C6774 XA2.XA4.MN0.G a_5960_47268# 0.155f
C6775 XA8.XA7.MP0.G a_19928_43748# 1.95e-19
C6776 XA2.XA1.XA5.MN2.G XA1.XA1.XA2.MP0.D 0.146f
C6777 VREF a_7328_45860# 0.0178f
C6778 XA2.XA4.MN0.D a_4808_45860# 2.24e-19
C6779 AVDD a_2288_40228# 0.464f
C6780 a_23600_47972# XA20.XA3a.MN0.D 0.00224f
C6781 XA2.XA11.MN1.G XA1.XA10.MP0.G 0.00598f
C6782 AVDD a_8480_52196# 0.00154f
C6783 DONE XA8.XA9.MN1.G 0.0317f
C6784 XA4.XA11.MP0.D a_11000_53252# 0.0494f
C6785 a_21080_53604# a_21080_53252# 0.0109f
C6786 a_17408_40580# a_17408_40228# 0.0109f
C6787 XA5.XA1.XA5.MN2.G a_12368_41284# 5.96e-19
C6788 XA6.XA4.MN0.G a_14888_44100# 0.0164f
C6789 XA7.XA6.MP0.G a_17408_42692# 5.5e-19
C6790 XA0.XA11.MN1.G a_9560_n18# 0.00214f
C6791 a_17408_46212# a_18560_46212# 0.00133f
C6792 XA3.XA6.MP0.G XA3.XA1.XA4.MP0.D 9.97e-19
C6793 XA6.XA3.MN0.G a_16040_45508# 0.0698f
C6794 XA6.XA9.MN1.G XA5.XA7.MP0.D 0.00108f
C6795 XA3.XA10.MP0.G a_8480_51492# 6.8e-20
C6796 AVDD a_19928_50084# 0.00154f
C6797 XA2.XA9.MN1.G a_4808_51844# 0.0164f
C6798 SARN a_23600_52196# 0.156f
C6799 CK_SAMPLE XA4.XA6.MP0.D 0.0276f
C6800 a_13808_1038# CK_SAMPLE_BSSW 5.11e-19
C6801 a_14960_1038# a_14960_686# 0.0109f
C6802 XB2.XA3.MN1.D a_13808_n18# 9.07e-19
C6803 XA20.XA3a.MN0.D a_22448_42340# 5.42e-19
C6804 a_11000_44452# a_12368_44452# 8.89e-19
C6805 XA6.XA6.MP0.G a_17408_39876# 1.28e-19
C6806 a_n232_44804# EN 9.82e-19
C6807 XA7.XA6.MP0.G a_13520_39876# 0.00296f
C6808 XA0.XA4.MN0.D a_920_40580# 9.14e-20
C6809 SARN li_14804_19176# 0.00103f
C6810 D<7> D<3> 9.11e-19
C6811 D<6> D<4> 0.568f
C6812 XA8.XA1.XA5.MN2.G a_16040_50788# 7.1e-20
C6813 XA7.XA1.XA5.MN2.G a_17408_50788# 7.1e-20
C6814 a_18560_51140# XA7.XA6.MN2.D 0.00176f
C6815 AVDD XA7.XA3.MN0.G 2.47f
C6816 XA6.XA9.MN1.G a_16040_49732# 0.0215f
C6817 XA2.XA9.MN1.G VREF 0.0732f
C6818 XA20.XA10.MN1.D a_22448_47972# 2.14e-19
C6819 XB2.XA4.MP0.D m3_16472_308# 0.106f
C6820 li_14804_20820# li_14804_20208# 0.00271f
C6821 XDAC2.XC128b<2>.XRES2.B XDAC2.XC128b<2>.XRES1A.B 0.0136f
C6822 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128a<1>.XRES4.B 0.00284f
C6823 XDAC1.XC128b<2>.XRES16.B li_9184_20208# 0.00117f
C6824 XA0.XA6.MP0.G XDAC2.XC32a<0>.XRES16.B 2.43e-19
C6825 EN XA3.XA1.XA4.MN0.D 3.17e-19
C6826 XA20.XA2a.MN0.D a_4808_40580# 0.00138f
C6827 XA1.XA1.XA2.MP0.D XA1.XA1.XA4.MN1.D 0.056f
C6828 XA5.XA1.XA2.MP0.D a_13520_43044# 0.0292f
C6829 XA5.XA1.XA5.MP0.D a_12368_43044# 0.00176f
C6830 a_11000_43396# a_12368_43396# 8.89e-19
C6831 XA1.XA4.MN0.D XDAC1.X16ab.XRES16.B 1.21e-19
C6832 XA7.XA6.MP0.G XA3.XA4.MN0.D 0.0254f
C6833 XA3.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.885f
C6834 XA3.XA6.MP0.G a_7328_49380# 0.0781f
C6835 XA8.XA6.MP0.G VREF 0.5f
C6836 XA20.XA3a.MN0.G a_22448_49732# 0.159f
C6837 AVDD a_23600_43748# 0.00154f
C6838 XA6.XA6.MP0.G XA6.XA4.MN0.D 0.76f
C6839 XA0.XA7.MP0.G a_920_47620# 0.00363f
C6840 SARP XB2.XA0.MP0.D 4.23e-19
C6841 a_22448_42340# a_23600_42340# 0.00133f
C6842 XA20.XA1.MN0.D a_22448_41988# 2.16e-19
C6843 XA5.XA1.XA5.MN2.G a_9848_44452# 1.86e-19
C6844 a_4808_48324# XA2.XA4.MN0.G 0.0677f
C6845 AVDD a_11000_41284# 0.361f
C6846 VREF a_5960_46916# 0.0536f
C6847 XA8.XA4.MN0.D a_21080_47268# 0.058f
C6848 XA20.XA3.MN6.D XA20.XA2a.MN0.D 0.431f
C6849 D<3> a_12368_45156# 6.68e-19
C6850 XA7.XA12.MP0.G XA8.XA12.MP0.G 0.00217f
C6851 AVDD a_5960_52900# 0.387f
C6852 a_19928_53956# a_19928_53604# 0.0109f
C6853 XA4.XA11.MN1.G a_7328_53604# 0.00979f
C6854 SARP li_9184_8736# 0.00103f
C6855 XA3.XA1.XA1.MN0.S a_8480_39876# 2.54e-19
C6856 XA8.XA1.XA1.MN0.S a_21080_40228# 0.0313f
C6857 a_9848_40932# a_11000_40932# 0.00133f
C6858 XA3.XA4.MN0.G a_7328_45156# 5.54e-19
C6859 XA3.XA3.MN0.G a_7328_46564# 0.155f
C6860 D<6> XA2.XA1.XA4.MP0.D 6.08e-19
C6861 XA7.XA1.XA5.MN2.G a_18560_42340# 0.00568f
C6862 XA8.XA1.XA5.MN2.G a_17408_42340# 0.00442f
C6863 XA0.XA7.MP0.G a_920_41988# 0.0719f
C6864 XA20.XA3.MN0.D a_23600_43748# 0.0765f
C6865 D<2> a_16040_42692# 7.76e-20
C6866 XA0.XA11.MN1.G XB2.XA2.MN0.G 0.0721f
C6867 XA5.XA10.MP0.G XA5.XA9.MN1.G 0.202f
C6868 a_3440_52548# XA1.XA9.MN1.G 0.0711f
C6869 a_14888_52548# a_16040_52548# 0.00133f
C6870 AVDD a_18560_50788# 0.00154f
C6871 CK_SAMPLE XA3.XA6.MP2.D 3.06e-19
C6872 SAR_IN XB2.XA0.MP0.D 0.115f
C6873 SAR_IP a_9560_1742# 0.0425f
C6874 XA4.XA6.MP0.G a_11000_40932# 4.24e-19
C6875 XA0.XA6.MP0.G a_920_40580# 5.5e-19
C6876 XA20.XA3a.MN0.D XA2.XA1.XA4.MN1.D 0.0124f
C6877 XA5.XA4.MN0.G a_12368_42692# 0.00224f
C6878 a_16040_53252# VREF 0.00292f
C6879 XA2.XA7.MP0.D a_4808_50788# 3.29e-19
C6880 XA6.XA9.MN1.G a_16040_50436# 7.76e-19
C6881 AVDD a_21080_47972# 0.356f
C6882 XA1.XA9.MN1.G XA1.XA6.MP0.G 0.0725f
C6883 XA3.XA1.XA5.MN2.G XA4.XA1.XA5.MN2.G 1.58f
C6884 a_21080_51492# XA8.XA7.MP0.G 0.0699f
C6885 a_9848_51492# a_9848_51140# 0.0109f
C6886 XA3.XA6.MP0.G XDAC2.X16ab.XRES8.B 0.00669f
C6887 XA0.XA1.XA2.MP0.D XA0.XA1.XA5.MP0.D 4.34e-19
C6888 XA8.XA1.XA5.MN1.D XA8.XA1.XA2.MP0.D 0.0102f
C6889 XA20.XA2a.MN0.D XA4.XA1.XA1.MP2.D 0.0102f
C6890 D<8> XA0.XA1.XA1.MN0.D 0.00135f
C6891 EN a_17408_43396# 0.162f
C6892 AVDD a_8480_44452# 0.00125f
C6893 D<0> a_21080_49732# 0.0109f
C6894 a_22448_50436# XA20.XA3a.MN0.G 0.0676f
C6895 D<3> XA5.XA4.MN0.D 0.203f
C6896 XA8.XA1.XA5.MN2.G a_16040_49028# 7.1e-20
C6897 XA7.XA1.XA5.MN2.G a_17408_49028# 7.1e-20
C6898 D<6> a_5960_49380# 0.00891f
C6899 D<1> XA0.XA4.MN0.D 0.0445f
C6900 D<2> XA2.XA4.MN0.D 5.62e-19
C6901 XA6.XA6.MP2.D VREF 5.13e-19
C6902 EN a_16040_40932# 0.00564f
C6903 D<8> li_14804_29616# 3.5e-20
C6904 XA6.XA1.XA2.MP0.D XA6.XA1.XA1.MN0.S 2.11e-19
C6905 a_14888_42692# XA6.XA1.XA4.MN0.D 0.00176f
C6906 SARN a_23600_44452# 0.0017f
C6907 XA20.XA3a.MN0.G a_23600_47620# 0.154f
C6908 XA20.XA3.MN6.D a_22448_47620# 0.00966f
C6909 XA5.XA6.MP0.G a_13520_47268# 1.38e-19
C6910 XA1.XA6.MP0.G a_3440_46916# 7.76e-20
C6911 a_21080_49028# a_22448_49028# 8.89e-19
C6912 XA5.XA1.XA5.MN2.G a_9848_45508# 2.31e-19
C6913 AVDD a_19928_42340# 0.00159f
C6914 VREF XA4.XA4.MN0.G 0.263f
C6915 XA8.XA4.MN0.D a_19928_48324# 0.0981f
C6916 XA2.XA4.MN0.D XA2.XA4.MN0.G 0.728f
C6917 AVDD XA6.XA12.MP0.G 0.709f
C6918 a_920_54308# XA0.XA12.MP0.D 0.00177f
C6919 a_920_41284# XA0.XA1.XA1.MP1.D 0.00176f
C6920 XA0.XA1.XA1.MP2.D a_920_40932# 0.00176f
C6921 XA5.XA1.XA1.MN0.S XA5.XA1.XA1.MP1.D 0.0615f
C6922 XA3.XA1.XA5.MN2.G XA2.XA1.XA4.MP1.D 0.00353f
C6923 a_16040_47268# a_17408_47268# 8.89e-19
C6924 XA2.XA4.MN0.D a_4808_44804# 9.25e-20
C6925 VREF a_7328_44804# 0.0691f
C6926 XA20.XA3a.MN0.D XA8.XA3.MN0.G 0.00428f
C6927 XA3.XA6.MP0.G XA3.XA1.XA5.MN1.D 7.41e-19
C6928 XA8.XA4.MN0.G XA20.XA2a.MN0.D 0.0122f
C6929 XA2.XA4.MN0.G a_5960_46212# 3.46e-19
C6930 AVDD XB1.M1.G 0.717f
C6931 XA8.XA10.MP0.D a_19928_52900# 0.128f
C6932 XA2.XA10.MP0.D XA2.XA10.MP0.G 0.194f
C6933 CK_SAMPLE a_19928_51844# 0.00102f
C6934 AVDD XA0.XA7.MP0.G 5.46f
C6935 a_14888_53604# XA6.XA9.MN1.G 7.36e-20
C6936 XA20.XA3a.MN0.D XA0.XA1.XA2.MP0.D 0.195f
C6937 XA5.XA6.MP0.G a_13520_41636# 7.76e-20
C6938 SARN XB1.XA0.MP0.D 4.8e-19
C6939 a_11000_45508# a_12368_45508# 8.89e-19
C6940 a_16040_45860# XA6.XA1.XA5.MN2.D 3.12e-20
C6941 XA7.XA4.MN0.G XA7.XA1.XA5.MP0.D 0.00138f
C6942 XA3.XA1.XA5.MN2.G a_4808_40228# 5.59e-19
C6943 XA6.XA3.MN0.G a_14888_44452# 0.0934f
C6944 XA5.XA9.MN1.G a_13520_51140# 0.0469f
C6945 AVDD a_18560_49028# 0.00154f
C6946 XA0.XA9.MN1.G XA0.XA6.MN2.D 0.126f
C6947 a_920_51844# a_920_51492# 0.0109f
C6948 a_8480_51844# XA3.XA8.MP0.D 0.0215f
C6949 CK_SAMPLE a_3440_49380# 0.00139f
C6950 XDAC1.XC0.XRES16.B XDAC1.XC0.XRES1A.B 0.454f
C6951 XDAC2.XC0.XRES16.B li_14804_30648# 0.00117f
C6952 a_5960_44100# a_5960_43748# 0.0109f
C6953 a_17408_44100# XA7.XA1.XA5.MP1.D 0.00176f
C6954 EN XA4.XA1.XA5.MN1.D 0.0157f
C6955 XA20.XA2a.MN0.D XA8.XA1.XA4.MP0.D 0.0269f
C6956 a_4808_44452# XA2.XA1.XA2.MP0.D 5.16e-20
C6957 XA0.XA6.MP2.G li_9184_24300# 3.5e-20
C6958 SARN XDAC2.XC1.XRES1B.B 3.59f
C6959 XA6.XA8.MP0.D VREF 7.83e-19
C6960 XA7.XA1.XA5.MN2.G a_17408_50084# 7.1e-20
C6961 XA8.XA1.XA5.MN2.G a_16040_50084# 7.1e-20
C6962 D<3> XA2.XA6.MP0.G 0.191f
C6963 D<2> XA1.XA6.MP0.G 0.0376f
C6964 a_21080_51140# XA8.XA6.MP0.G 6.76e-20
C6965 D<1> XA0.XA6.MP0.G 0.173f
C6966 XA8.XA6.MN2.D a_19928_50436# 0.00176f
C6967 a_8480_50788# a_8480_50436# 0.0109f
C6968 D<4> XA3.XA6.MP0.G 0.0877f
C6969 AVDD a_8480_45508# 0.00131f
C6970 D<0> a_21080_50436# 0.0879f
C6971 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES8.B 0.0228f
C6972 XDAC1.XC128a<1>.XRES16.B XDAC1.XC32a<0>.XRES16.B 0.0114f
C6973 li_9184_15696# li_9184_15084# 0.00271f
C6974 XA2.XA1.XA4.MN1.D XA2.XA1.XA4.MP1.D 0.00918f
C6975 XA0.XA4.MN0.D XDAC1.XC32a<0>.XRES16.B 2.43e-19
C6976 EN a_22448_41636# 5.7e-20
C6977 AVDD XA1.XA1.XA4.MP1.D 0.0913f
C6978 XA6.XA1.XA5.MN2.G XA6.XA3.MN0.G 5.78e-19
C6979 XA2.XA1.XA5.MN2.G a_920_46564# 7.1e-20
C6980 XA0.XA7.MP0.G a_2288_46564# 7.1e-20
C6981 XA20.XA10.MN1.D a_23600_43748# 0.00405f
C6982 VREF a_16040_49380# 0.0171f
C6983 XA4.XA4.MN0.D a_11000_49380# 0.154f
C6984 a_21080_49732# a_21080_49380# 0.0109f
C6985 SARN a_23600_45508# 0.0017f
C6986 XA5.XA6.MP0.G a_12368_48324# 0.00417f
C6987 XA20.XA3a.MN0.G a_22448_48676# 0.0268f
C6988 a_16040_41636# a_17408_41636# 8.89e-19
C6989 SARP XDAC1.XC64b<1>.XRES4.B 13.9f
C6990 XA2.XA4.MN0.G a_4808_47268# 0.157f
C6991 XA8.XA1.XA5.MN2.G a_19928_43748# 0.0732f
C6992 XA0.XA7.MP0.G XA1.XA1.XA2.MP0.D 0.126f
C6993 VREF a_5960_45860# 0.0178f
C6994 AVDD a_920_40228# 0.467f
C6995 a_22448_47972# XA20.XA3a.MN0.D 0.00239f
C6996 AVDD a_7328_52196# 0.37f
C6997 XA6.XA11.MN1.G a_14888_52900# 7.39e-19
C6998 XA5.XA12.MP0.G a_13520_52900# 0.00258f
C6999 a_920_53252# a_2288_53252# 8.89e-19
C7000 a_3440_40228# a_4808_40228# 8.89e-19
C7001 XA5.XA1.XA5.MN2.G a_11000_41284# 0.0175f
C7002 XA6.XA4.MN0.G a_13520_44100# 2.84e-19
C7003 XA5.XA4.MN0.G a_14888_44100# 2.84e-19
C7004 XA0.XA4.MN0.D a_920_43044# 9.14e-20
C7005 a_4808_46212# a_4808_45860# 0.0109f
C7006 XA6.XA3.MN0.G a_14888_45508# 0.104f
C7007 AVDD a_18560_50084# 0.00144f
C7008 CK_SAMPLE XA4.XA6.MN0.D 0.0659f
C7009 XA2.XA9.MN1.G a_3440_51844# 2.2e-19
C7010 XA5.XA9.MN0.D XA5.XA7.MP0.D 0.00986f
C7011 a_9848_52196# a_11000_52196# 0.00133f
C7012 XA5.XA9.MN1.G XA6.XA7.MP0.D 0.00108f
C7013 a_7328_52900# XA4.XA1.XA5.MN2.G 1.06e-19
C7014 a_9560_686# a_11000_686# 8e-19
C7015 XA20.XA3a.MN0.D a_21080_42340# 8.09e-19
C7016 XA20.XA2a.MN0.D a_4808_43044# 1.43e-19
C7017 XA3.XA1.XA5.MN2.D a_8480_43748# 0.00224f
C7018 XA6.XA6.MP0.G a_16040_39876# 0.00207f
C7019 XA2.XA4.MN0.G a_4808_41636# 6.69e-20
C7020 SARP a_23600_44452# 0.154f
C7021 XA7.XA6.MP0.G a_12368_39876# 0.00332f
C7022 XA0.XA4.MN0.D a_n232_40580# 9.25e-20
C7023 a_5960_51140# a_5960_50788# 0.0109f
C7024 XA7.XA1.XA5.MN2.G a_16040_50788# 0.00548f
C7025 AVDD XA6.XA3.MN0.G 2.47f
C7026 XA1.XA9.MN1.G XA1.XA4.MN0.D 0.00938f
C7027 XA6.XA9.MN1.G a_14888_49732# 0.00119f
C7028 XA2.XA7.MP0.D a_4808_50084# 7.44e-20
C7029 XB2.XA4.MP0.D m3_26048_1188# 0.0273f
C7030 XB1.XA3.MN1.D m3_n1960_132# 0.0634f
C7031 EN XA3.XA1.XA4.MP0.D 0.0386f
C7032 XA20.XA2a.MN0.D a_3440_40580# 0.00123f
C7033 XA5.XA1.XA2.MP0.D a_12368_43044# 3.59e-19
C7034 XA1.XA1.XA2.MP0.D XA1.XA1.XA4.MP1.D 4.34e-19
C7035 a_21080_50084# a_22448_50084# 8.89e-19
C7036 a_8480_50084# a_8480_49732# 0.0109f
C7037 XA8.XA1.XA5.MN2.G a_17408_47972# 0.00363f
C7038 D<0> a_21080_48676# 0.00918f
C7039 XA2.XA1.XA5.MN2.G XA20.XA3a.MN0.D 0.963f
C7040 D<4> a_11000_48324# 0.0164f
C7041 AVDD a_22448_43748# 0.491f
C7042 SARP XB1.XA0.MP0.D 0.00704f
C7043 a_9848_42340# a_9848_41988# 0.0109f
C7044 D<8> XDAC2.XC128a<1>.XRES1B.B 0.00406f
C7045 XA4.XA1.XA5.MN2.G a_9848_44452# 5.11e-19
C7046 a_14888_48324# a_16040_48324# 0.00133f
C7047 AVDD a_9848_41284# 0.00125f
C7048 XA1.XA4.MN0.D a_3440_46916# 0.00456f
C7049 XA8.XA4.MN0.D a_19928_47268# 0.0963f
C7050 XA5.XA6.MP0.G a_13520_46212# 4.4e-19
C7051 XA20.XA3a.MN0.G XA20.XA2a.MN0.D 0.222f
C7052 XA20.XA3.MN6.D a_23600_46564# 0.0665f
C7053 XA1.XA6.MP0.G a_3440_45860# 7.76e-20
C7054 AVDD a_4808_52900# 0.00166f
C7055 XA20.XA12.MP0.D XA20.XA9.MP0.D 2.14e-19
C7056 XA20.XA12.MP0.G XA8.XA10.MP0.D 0.00171f
C7057 XA3.XA11.MN1.G a_8480_53604# 0.0726f
C7058 XA4.XA11.MN1.G a_5960_53604# 9.49e-20
C7059 XA8.XA11.MN1.G XA8.XA12.MP0.G 0.214f
C7060 XA3.XA1.XA1.MN0.S a_7328_39876# 2.54e-19
C7061 XA8.XA1.XA1.MN0.S a_19928_40228# 0.0215f
C7062 XA3.XA1.XA1.MN0.D a_8480_40580# 0.035f
C7063 XA8.XA1.XA1.MP1.D a_21080_40932# 0.0465f
C7064 a_17408_46916# a_17408_46564# 0.0109f
C7065 D<6> XA2.XA1.XA4.MN0.D 0.00144f
C7066 XA7.XA1.XA5.MN2.G a_17408_42340# 1.97e-19
C7067 XA0.XA7.MP0.G a_n232_41988# 0.0684f
C7068 XA4.XA6.MP0.G a_11000_43396# 5.5e-19
C7069 VREF XA7.XA1.XA5.MP1.D 0.00623f
C7070 D<2> a_14888_42692# 6.49e-19
C7071 XA0.XA6.MP0.G a_920_43044# 5.5e-19
C7072 a_2288_52548# XA1.XA9.MN1.G 0.0674f
C7073 AVDD a_17408_50788# 0.363f
C7074 CK_SAMPLE D<5> 0.0524f
C7075 XB2.XA1.MN0.D XB2.XA0.MP0.D 0.0115f
C7076 SAR_IP a_8408_1742# 0.0215f
C7077 a_14960_2446# XB2.XA4.MP0.D 0.00977f
C7078 XB2.XA1.MP0.D a_14960_2094# 2.01e-19
C7079 a_11000_2446# a_11000_2094# 0.0109f
C7080 a_14960_3150# XB2.XA3.MN1.D 0.00238f
C7081 XB1.XA1.MN0.D a_9560_1742# 1.71e-19
C7082 XA4.XA6.MP0.G a_9848_40932# 3.97e-20
C7083 XA0.XA6.MP0.G a_n232_40580# 7.76e-20
C7084 SARN li_14804_29616# 0.00103f
C7085 XA20.XA3a.MN0.D XA1.XA1.XA4.MN1.D 0.0124f
C7086 XA6.XA1.XA5.MN2.D a_16040_44804# 0.156f
C7087 a_5960_45156# a_5960_44804# 0.0109f
C7088 XA20.XA2a.MN0.D a_n232_43748# 4.48e-20
C7089 D<3> a_14888_39876# 1.26e-19
C7090 a_18560_45156# a_19928_45156# 8.89e-19
C7091 XA6.XA9.MN1.G a_14888_50436# 0.01f
C7092 AVDD a_19928_47972# 0.00159f
C7093 XA8.XA7.MP0.D D<0> 1.69e-19
C7094 a_19928_51492# XA8.XA7.MP0.G 0.0674f
C7095 XDAC2.XC64b<1>.XRES16.B XDAC2.X16ab.XRES16.B 0.0114f
C7096 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES8.B 0.0228f
C7097 li_14804_26136# li_14804_25524# 0.00271f
C7098 a_9848_43748# XA4.XA1.XA5.MN0.D 0.00176f
C7099 XA3.XA1.XA5.MP1.D a_7328_43396# 0.00176f
C7100 XA0.XA1.XA2.MP0.D XA0.XA1.XA5.MN0.D 0.056f
C7101 XA20.XA2a.MN0.D XA4.XA1.XA1.MN0.S 0.137f
C7102 EN a_16040_43396# 0.162f
C7103 XA0.XA6.MP0.G XDAC2.X16ab.XRES16.B 2.4e-19
C7104 AVDD a_7328_44452# 0.357f
C7105 XA1.XA6.MP0.G XA7.XA6.MP0.G 0.0649f
C7106 D<0> a_19928_49732# 7.01e-19
C7107 XA7.XA1.XA5.MN2.G a_16040_49028# 0.00363f
C7108 D<6> a_4808_49380# 5.91e-19
C7109 XA2.XA6.MP0.G XA6.XA6.MP0.G 0.047f
C7110 XA3.XA6.MP0.G XA5.XA6.MP0.G 0.059f
C7111 D<2> XA1.XA4.MN0.D 0.0331f
C7112 a_8480_50436# a_8480_50084# 0.0109f
C7113 XDAC2.XC64a<0>.XRES2.B XDAC2.XC64a<0>.XRES16.B 0.457f
C7114 XDAC2.XC64a<0>.XRES8.B XDAC2.XC64a<0>.XRES1A.B 0.0228f
C7115 XA2.XA1.XA2.MP0.D a_5960_41284# 1.07e-19
C7116 XA5.XA1.XA4.MN1.D a_13520_42340# 0.00176f
C7117 a_2288_42692# a_2288_42340# 0.0109f
C7118 XA1.XA3.MN0.G XDAC2.XC64b<1>.XRES1B.B 0.00405f
C7119 XA20.XA3a.MN0.G a_22448_47620# 0.181f
C7120 XA5.XA6.MP0.G a_12368_47268# 5.95e-19
C7121 XA1.XA6.MP0.G a_2288_46916# 5.5e-19
C7122 a_8480_49028# a_8480_48676# 0.0109f
C7123 XA4.XA1.XA5.MN2.G a_9848_45508# 9.01e-20
C7124 AVDD a_18560_42340# 0.00125f
C7125 VREF XA3.XA4.MN0.G 0.263f
C7126 XA1.XA4.MN0.D XA2.XA4.MN0.G 3.16e-20
C7127 XA2.XA4.MN0.D XA1.XA4.MN0.G 3.16e-20
C7128 AVDD XA7.XA11.MN1.G 1.89f
C7129 a_n232_54308# XA0.XA12.MP0.D 2.54e-19
C7130 a_12368_54308# a_12368_53956# 0.0109f
C7131 SARP li_9184_19176# 0.00103f
C7132 a_12368_41284# a_13520_41284# 0.00133f
C7133 XA0.XA1.XA1.MN0.S a_920_40932# 0.0271f
C7134 D<1> XA7.XA1.XA5.MN0.D 0.00188f
C7135 XA3.XA1.XA5.MN2.G XA2.XA1.XA4.MN1.D 7.2e-19
C7136 a_3440_47268# a_3440_46916# 0.0109f
C7137 XA8.XA7.MP0.G a_22448_43044# 0.00113f
C7138 VREF a_5960_44804# 0.0691f
C7139 XA2.XA1.XA5.MN2.G XA2.XA1.XA4.MP1.D 7.44e-19
C7140 XA7.XA6.MP0.G a_18560_44100# 7.76e-20
C7141 XA20.XA3a.MN0.D XA7.XA3.MN0.G 7.15e-20
C7142 XA3.XA6.MP0.G XA3.XA1.XA5.MP1.D 0.00121f
C7143 XA7.XA4.MN0.G XA20.XA2a.MN0.D 0.00833f
C7144 XA2.XA4.MN0.G a_4808_46212# 0.0149f
C7145 AVDD a_14960_2446# 0.406f
C7146 a_7328_52900# a_8480_52900# 0.00133f
C7147 CK_SAMPLE a_18560_51844# 2.08e-19
C7148 AVDD a_23600_51492# 0.00183f
C7149 XA2.XA11.MN1.G XA1.XA7.MP0.D 4.87e-19
C7150 a_22448_39876# a_23600_39876# 0.00133f
C7151 XA5.XA6.MP0.G a_12368_41636# 5.5e-19
C7152 XA1.XA6.MP0.G XA1.XA1.XA1.MN0.S 0.0123f
C7153 a_23600_45860# a_23600_45508# 0.0109f
C7154 XA0.XA4.MN0.G a_920_43396# 8.07e-19
C7155 XA7.XA4.MN0.G XA7.XA1.XA2.MP0.D 0.206f
C7156 XA8.XA7.MP0.G a_21080_40580# 0.0436f
C7157 XA2.XA1.XA5.MN2.G a_4808_40228# 0.0709f
C7158 D<5> a_8480_40932# 5.26e-19
C7159 XA5.XA9.MN1.G a_12368_51140# 0.0222f
C7160 AVDD a_17408_49028# 0.356f
C7161 XA0.XA9.MN1.G XA0.XA6.MP2.G 0.0378f
C7162 a_7328_51844# XA3.XA8.MP0.D 0.0215f
C7163 a_17408_51844# a_18560_51844# 0.00133f
C7164 XA3.XA7.MP0.D a_8480_51492# 0.126f
C7165 CK_SAMPLE a_2288_49380# 7.89e-19
C7166 a_12368_53956# VREF 0.00396f
C7167 D<5> XDAC1.X16ab.XRES4.B 0.00405f
C7168 EN XA3.XA1.XA5.MN1.D 0.0157f
C7169 XA20.XA2a.MN0.D XA8.XA1.XA4.MN0.D 0.0397f
C7170 XA4.XA1.XA5.MN2.D a_11000_43044# 1.88e-19
C7171 a_14888_44804# XA6.XA1.XA2.MP0.D 2.6e-20
C7172 XA2.XA3.MN0.G a_4808_41988# 0.00335f
C7173 XA5.XA8.MP0.D VREF 7.83e-19
C7174 D<5> XA3.XA6.MN0.D 0.00148f
C7175 AVDD a_7328_45508# 0.359f
C7176 a_19928_50788# a_21080_50788# 0.00133f
C7177 D<0> a_19928_50436# 5.7e-19
C7178 XA7.XA1.XA5.MN2.G a_16040_50084# 0.00366f
C7179 a_5960_43044# a_5960_42692# 0.0109f
C7180 a_17408_43044# XA7.XA1.XA4.MP1.D 0.00176f
C7181 EN a_21080_41636# 0.00643f
C7182 XA20.XA10.MN1.D a_22448_43748# 1.97e-19
C7183 VREF a_14888_49380# 8.08e-19
C7184 XA4.XA4.MN0.D a_9848_49380# 0.155f
C7185 AVDD XA0.XA1.XA4.MP1.D 0.0913f
C7186 D<4> a_11000_47268# 0.0148f
C7187 XA6.XA1.XA5.MN2.G XA5.XA3.MN0.G 0.106f
C7188 XA0.XA6.MP2.G a_920_46916# 0.0185f
C7189 XA0.XA7.MP0.G a_920_46564# 0.00363f
C7190 a_920_49380# a_2288_49380# 8.89e-19
C7191 D<0> a_21080_47620# 0.0147f
C7192 XA1.XA6.MP0.G XA1.XA4.MN0.G 0.0407f
C7193 XA20.XA3.MN6.D XA8.XA1.XA5.MN2.D 0.00869f
C7194 XA1.XA6.MP0.G a_3440_44804# 7.76e-20
C7195 a_9848_47972# a_9848_47620# 0.0109f
C7196 XA8.XA4.MN0.G a_21080_47620# 0.155f
C7197 XA7.XA1.XA5.MN2.G a_19928_43748# 7.1e-20
C7198 XA8.XA1.XA5.MN2.G a_18560_43748# 2.66e-19
C7199 XA0.XA7.MP0.G XA0.XA1.XA5.MP0.D 0.00353f
C7200 XA8.XA4.MN0.D a_19928_46212# 1.1e-19
C7201 XA1.XA4.MN0.D a_3440_45860# 2.23e-19
C7202 VREF a_4808_45860# 1.19e-19
C7203 AVDD a_n232_40228# 0.00131f
C7204 a_22448_47972# a_23600_47972# 0.00133f
C7205 D<6> XA2.XA1.XA5.MP1.D 7.42e-19
C7206 D<4> EN 0.0683f
C7207 XA6.XA11.MN1.G a_13520_52900# 0.00295f
C7208 XA5.XA12.MP0.G a_12368_52900# 1.28e-19
C7209 XA0.XA12.MP0.D XA1.XA10.MP0.G 0.0119f
C7210 a_9848_53604# XA4.XA10.MP0.D 1.17e-19
C7211 a_19928_53604# a_19928_53252# 0.0109f
C7212 AVDD a_5960_52196# 0.37f
C7213 a_16040_40580# a_16040_40228# 0.0109f
C7214 D<4> a_11000_41636# 7.76e-20
C7215 XA5.XA1.XA5.MN2.G a_9848_41284# 0.00527f
C7216 XA5.XA4.MN0.G a_13520_44100# 0.0164f
C7217 XA0.XA4.MN0.D a_n232_43044# 9.25e-20
C7218 XA20.XA3a.MN0.D a_8480_44452# 2.59e-20
C7219 a_16040_46212# a_17408_46212# 8.89e-19
C7220 XA1.XA9.MN1.G a_4808_51844# 2.2e-19
C7221 XA1.XA9.MN0.D a_3440_51844# 0.00176f
C7222 AVDD a_17408_50084# 0.358f
C7223 CK_SAMPLE XA4.XA6.MP0.G 0.046f
C7224 XA5.XA9.MN1.G XA5.XA7.MP0.D 0.274f
C7225 a_13808_1038# a_13808_686# 0.0109f
C7226 XA20.XA3a.MN0.D a_19928_42340# 0.0059f
C7227 a_9848_44452# a_11000_44452# 0.00133f
C7228 XA20.XA2a.MN0.D a_3440_43044# 1.43e-19
C7229 XA3.XA1.XA5.MN2.D a_7328_43748# 0.00388f
C7230 XA6.XA6.MP0.G a_14888_39876# 8.17e-19
C7231 XA8.XA4.MN0.G a_21080_41988# 5.1e-20
C7232 XA20.XA2.MN1.D a_23600_44100# 0.0605f
C7233 a_23600_44804# a_23600_44452# 0.0109f
C7234 SARN XDAC2.XC128a<1>.XRES1B.B 3.59f
C7235 XA7.XA1.XA5.MN2.G a_14888_50788# 1.87e-19
C7236 a_17408_51140# XA7.XA6.MP2.D 0.00176f
C7237 AVDD XA5.XA3.MN0.G 2.47f
C7238 XA1.XA9.MN1.G VREF 0.0732f
C7239 XB2.XA4.MP0.D m3_25976_1188# 0.0137f
C7240 XB1.XA3.MN1.D m3_n2104_132# 0.17f
C7241 li_9184_20820# li_9184_20208# 0.00271f
C7242 XDAC1.XC128b<2>.XRES2.B XDAC1.XC128b<2>.XRES1A.B 0.0136f
C7243 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128a<1>.XRES4.B 0.00284f
C7244 EN XA2.XA1.XA4.MP0.D 0.0386f
C7245 XA0.XA6.MP0.G li_14804_13860# 1.85e-20
C7246 a_9848_43396# a_11000_43396# 0.00133f
C7247 XA3.XA3.MN0.G a_9848_40228# 9.08e-19
C7248 XA0.XA4.MN0.D XDAC1.X16ab.XRES16.B 2.4e-19
C7249 XA7.XA6.MP0.D VREF 0.0115f
C7250 XA7.XA1.XA5.MN2.G a_17408_47972# 7.1e-20
C7251 XA8.XA1.XA5.MN2.G a_16040_47972# 7.1e-20
C7252 D<0> a_19928_48676# 3.48e-19
C7253 XA0.XA7.MP0.G XA20.XA3a.MN0.D 0.885f
C7254 XA8.XA6.MP0.D a_21080_49732# 0.00176f
C7255 XA0.XA6.MP2.G XA0.XA4.MN0.G 0.259f
C7256 D<4> a_9848_48324# 6.53e-19
C7257 AVDD a_21080_43748# 0.357f
C7258 a_21080_42340# a_22448_42340# 8.89e-19
C7259 XA8.XA1.XA4.MP0.D a_21080_41988# 0.00176f
C7260 XA4.XA1.XA5.MN2.G a_8480_44452# 1.86e-19
C7261 XA8.XA4.MN0.D a_18560_47268# 4.76e-20
C7262 XA7.XA4.MN0.D a_19928_47268# 4.76e-20
C7263 XA1.XA4.MN0.D a_2288_46916# 0.00254f
C7264 AVDD a_8480_41284# 0.00125f
C7265 XA5.XA6.MP0.G a_12368_46212# 5.5e-19
C7266 XA20.XA3.MN6.D a_22448_46564# 0.0781f
C7267 XA20.XA3a.MN0.G a_23600_46564# 0.0677f
C7268 D<0> XA8.XA1.XA5.MN2.D 0.00547f
C7269 XA1.XA6.MP0.G a_2288_45860# 5.5e-19
C7270 a_3440_48324# XA1.XA4.MN0.G 0.0661f
C7271 a_19928_48676# XA8.XA4.MN0.G 1.34e-19
C7272 AVDD a_3440_52900# 0.00166f
C7273 a_18560_53956# a_18560_53604# 0.0109f
C7274 XA2.XA12.MP0.G a_5960_53604# 0.0893f
C7275 XA3.XA11.MN1.G a_7328_53604# 0.073f
C7276 XA8.XA11.MN1.G XA7.XA12.MP0.G 0.391f
C7277 SARP XDAC1.XC1.XRES1B.B 3.59f
C7278 XA3.XA1.XA1.MN0.D a_7328_40580# 8.3e-19
C7279 XA8.XA1.XA1.MN0.D a_21080_40932# 8.29e-20
C7280 a_8480_40932# a_9848_40932# 8.89e-19
C7281 XA8.XA4.MN0.G XA8.XA1.XA5.MN2.D 0.135f
C7282 XA2.XA4.MN0.G a_5960_45156# 5.54e-19
C7283 XA2.XA3.MN0.G a_5960_46564# 0.155f
C7284 XA7.XA1.XA5.MN2.G a_16040_42340# 0.00442f
C7285 XA4.XA6.MP0.G a_9848_43396# 7.76e-20
C7286 VREF XA6.XA1.XA5.MP1.D 0.00623f
C7287 XA0.XA6.MP0.G a_n232_43044# 7.76e-20
C7288 XA0.XA11.MN1.G a_13808_3502# 0.0379f
C7289 SARN a_23600_41284# 5.16e-19
C7290 XA4.XA10.MP0.G XA4.XA9.MN0.D 0.106f
C7291 a_13520_52548# a_14888_52548# 8.89e-19
C7292 XA20.XA10.MN1.D a_23600_51492# 0.0046f
C7293 CK_SAMPLE XA2.XA6.MP2.D 3.06e-19
C7294 AVDD a_16040_50788# 0.363f
C7295 XB1.M1.G XB2.M1.G 0.0182f
C7296 XB1.XA4.MP0.D XB1.XA4.MN0.D 0.00106f
C7297 XB2.XA1.MP0.D a_13808_2094# 0.0722f
C7298 a_8408_2798# XB1.XA3.MN1.D 3.55e-19
C7299 XB1.XA1.MP0.D a_9560_1742# 8.33e-19
C7300 XA1.XA4.MN0.D XA1.XA1.XA1.MN0.S 0.0145f
C7301 XA20.XA3a.MN0.D XA1.XA1.XA4.MP1.D 0.0124f
C7302 XA6.XA1.XA5.MN2.D a_14888_44804# 0.153f
C7303 D<3> a_13520_39876# 0.00212f
C7304 XA4.XA4.MN0.G a_11000_42692# 0.00224f
C7305 XA2.XA3.MN0.G XA2.XA1.XA2.MP0.D 0.0351f
C7306 AVDD a_18560_47972# 0.00125f
C7307 a_8480_51492# a_8480_51140# 0.0109f
C7308 XA2.XA1.XA5.MN2.G XA3.XA1.XA5.MN2.G 0.0255f
C7309 XA1.XA7.MP0.D a_3440_50788# 3.29e-19
C7310 a_9848_43748# XA4.XA1.XA2.MP0.D 0.0702f
C7311 XA7.XA1.XA5.MN1.D XA7.XA1.XA5.MN0.D 0.0488f
C7312 XA20.XA2a.MN0.D XA3.XA1.XA1.MP2.D 0.0102f
C7313 EN a_14888_43396# 0.00238f
C7314 AVDD a_5960_44452# 0.357f
C7315 a_21080_50436# XA8.XA6.MP0.D 0.00176f
C7316 D<3> XA3.XA4.MN0.D 0.0297f
C7317 D<2> VREF 1.3f
C7318 a_13520_42692# XA5.XA1.XA4.MN0.D 0.00176f
C7319 D<8> XDAC2.XC64b<1>.XRES1B.B 4.06e-21
C7320 a_19928_49028# a_21080_49028# 0.00133f
C7321 XA0.XA6.MP2.G a_920_45860# 0.0774f
C7322 XA4.XA1.XA5.MN2.G a_8480_45508# 2.31e-19
C7323 D<4> a_11000_46212# 0.0202f
C7324 AVDD a_17408_42340# 0.361f
C7325 VREF XA2.XA4.MN0.G 0.263f
C7326 XA7.XA4.MN0.D a_18560_48324# 0.0997f
C7327 XA1.XA4.MN0.D XA1.XA4.MN0.G 0.728f
C7328 AVDD XA5.XA12.MP0.G 0.706f
C7329 a_n232_41284# XA0.XA1.XA1.MN0.D 0.00224f
C7330 XA4.XA1.XA1.MP2.D XA4.XA1.XA1.MP1.D 0.0488f
C7331 D<1> XA7.XA1.XA5.MP0.D 7.43e-19
C7332 a_14888_47268# a_16040_47268# 0.00133f
C7333 XA8.XA7.MP0.G a_21080_43044# 0.00551f
C7334 VREF a_4808_44804# 7.12e-19
C7335 XA1.XA4.MN0.D a_3440_44804# 9.24e-20
C7336 XA2.XA1.XA5.MN2.G XA2.XA1.XA4.MN1.D 0.0131f
C7337 D<5> a_8480_43396# 6.49e-19
C7338 XA7.XA6.MP0.G a_17408_44100# 5.5e-19
C7339 XA20.XA3a.MN0.D XA6.XA3.MN0.G 7.15e-20
C7340 XA5.XA6.MP0.G EN 0.071f
C7341 XA6.XA4.MN0.G XA20.XA2a.MN0.D 0.00823f
C7342 XA1.XA4.MN0.G a_4808_46212# 2.2e-19
C7343 XA2.XA4.MN0.G a_3440_46212# 2.2e-19
C7344 AVDD a_13808_2446# 0.00166f
C7345 AVDD a_22448_51492# 0.568f
C7346 XA1.XA10.MP0.D XA1.XA10.MP0.G 0.194f
C7347 XA7.XA10.MP0.D a_18560_52900# 0.13f
C7348 XA20.XA3a.MN0.D a_22448_43748# 0.00726f
C7349 a_9848_45508# a_11000_45508# 0.00133f
C7350 XA0.XA4.MN0.G a_n232_43396# 0.0104f
C7351 XA5.XA3.MN0.G a_13520_44452# 0.0934f
C7352 XA8.XA7.MP0.G a_19928_40580# 1.39e-19
C7353 XA8.XA1.XA5.MN2.G a_21080_40580# 6.02e-19
C7354 XA2.XA1.XA5.MN2.G a_3440_40228# 1.34e-19
C7355 XA0.XA7.MP0.G a_4808_40228# 4.72e-19
C7356 D<5> a_7328_40932# 4.18e-20
C7357 SARN a_13808_2094# 0.00112f
C7358 AVDD a_16040_49028# 0.356f
C7359 a_n232_51844# a_n232_51492# 0.0109f
C7360 XA3.XA7.MP0.D a_7328_51492# 0.0877f
C7361 CK_SAMPLE a_920_49380# 7.89e-19
C7362 a_11000_53956# VREF 0.00366f
C7363 a_7328_52196# XA4.XA1.XA5.MN2.G 3.39e-19
C7364 XDAC2.XC0.XRES4.B XDAC2.XC64b<1>.XRES4.B 0.00284f
C7365 li_14804_31260# li_14804_30648# 0.00271f
C7366 XDAC2.XC0.XRES2.B XDAC2.XC0.XRES1A.B 0.0136f
C7367 XDAC1.XC0.XRES16.B li_9184_30648# 0.00117f
C7368 a_4808_44100# a_4808_43748# 0.0109f
C7369 a_16040_44100# XA6.XA1.XA5.MP1.D 0.00176f
C7370 EN XA3.XA1.XA5.MP1.D 0.0543f
C7371 XA1.XA1.XA5.MP1.D XA1.XA1.XA5.MN1.D 0.00918f
C7372 XA20.XA3a.MN0.D a_9848_41284# 0.00649f
C7373 XA20.XA2a.MN0.D XA7.XA1.XA4.MN0.D 0.0409f
C7374 XA4.XA1.XA5.MN2.D a_9848_43044# 5.1e-20
C7375 XA0.XA6.MP2.G XDAC1.X16ab.XRES2.B 4.06e-21
C7376 SARN li_14804_9156# 0.00103f
C7377 XA1.XA3.MN0.G a_4808_41988# 4.4e-20
C7378 XA2.XA3.MN0.G a_3440_41988# 4.21e-19
C7379 XA4.XA8.MP0.D VREF 7.83e-19
C7380 a_7328_50788# a_7328_50436# 0.0109f
C7381 AVDD a_5960_45508# 0.359f
C7382 D<5> XA3.XA6.MP0.D 0.0323f
C7383 XDAC2.XC32a<0>.XRES1B.B XDAC2.XC32a<0>.XRES4.B 0.428f
C7384 XA7.XA1.XA2.MP0.D XA7.XA1.XA4.MN0.D 0.056f
C7385 SARP a_23600_41284# 0.16f
C7386 XA0.XA4.MN0.D li_9184_13860# 1.85e-20
C7387 EN a_19928_41636# 1.25e-19
C7388 VREF a_13520_49380# 8.08e-19
C7389 a_19928_49732# a_19928_49380# 0.0109f
C7390 AVDD XA0.XA1.XA4.MN1.D 0.00889f
C7391 D<4> a_9848_47268# 3.18e-19
C7392 XA6.XA1.XA5.MN2.G XA4.XA3.MN0.G 6.95e-19
C7393 XA5.XA1.XA5.MN2.G XA5.XA3.MN0.G 0.00127f
C7394 XA0.XA6.MP2.G a_n232_46916# 0.00249f
C7395 D<0> a_19928_47620# 5.21e-19
C7396 a_16040_41988# XA6.XA1.XA1.MN0.S 3.8e-19
C7397 a_14888_41636# a_16040_41636# 0.00133f
C7398 a_3440_41636# XA1.XA1.XA1.MN0.S 0.0658f
C7399 a_2288_41636# XA1.XA1.XA1.MP2.D 0.00176f
C7400 SARP li_9184_29616# 0.00103f
C7401 XA1.XA6.MP0.G a_2288_44804# 5.5e-19
C7402 D<2> a_16040_44100# 7.76e-20
C7403 XA1.XA4.MN0.G a_3440_47268# 0.157f
C7404 XA8.XA4.MN0.G a_19928_47620# 0.154f
C7405 XA8.XA1.XA5.MN2.G a_17408_43748# 0.00442f
C7406 XA7.XA1.XA5.MN2.G a_18560_43748# 0.0749f
C7407 XA0.XA7.MP0.G XA0.XA1.XA5.MN0.D 7.2e-19
C7408 XA1.XA4.MN0.D a_2288_45860# 9.15e-20
C7409 VREF a_3440_45860# 1.19e-19
C7410 AVDD a_23600_40580# 0.00181f
C7411 D<6> XA2.XA1.XA5.MN1.D 0.00185f
C7412 XA5.XA6.MP0.G a_13520_45156# 7.76e-20
C7413 XA6.XA11.MN1.G a_12368_52900# 1.34e-19
C7414 a_n232_53252# a_920_53252# 0.00133f
C7415 XA0.XA12.MP0.D XA0.XA10.MP0.G 0.0024f
C7416 AVDD a_4808_52196# 0.00154f
C7417 a_2288_40228# a_3440_40228# 0.00133f
C7418 D<4> a_9848_41636# 6.49e-19
C7419 XA4.XA1.XA5.MN2.G a_9848_41284# 0.0044f
C7420 XA0.XA6.MP2.G XA0.XA1.XA1.MN0.S 0.0149f
C7421 XA5.XA4.MN0.G a_12368_44100# 6.11e-19
C7422 XA0.XA11.MN1.G a_13808_334# 0.00214f
C7423 a_3440_46212# a_3440_45860# 0.0109f
C7424 XA5.XA3.MN0.G a_13520_45508# 0.106f
C7425 XA1.XA9.MN1.G a_3440_51844# 0.0164f
C7426 AVDD a_16040_50084# 0.358f
C7427 CK_SAMPLE XA3.XA6.MN0.D 0.0676f
C7428 a_8480_52196# a_9848_52196# 8.89e-19
C7429 XA20.XA9.MP0.D XA8.XA7.MP0.G 0.0216f
C7430 a_5960_52900# XA3.XA1.XA5.MN2.G 1.06e-19
C7431 a_9560_1038# CK_SAMPLE_BSSW 5.11e-19
C7432 a_8408_686# a_9560_686# 0.00133f
C7433 XA20.XA3a.MN0.D a_18560_42340# 0.00552f
C7434 XA6.XA6.MP0.G a_13520_39876# 7.4e-19
C7435 XA8.XA4.MN0.G a_19928_41988# 1.74e-19
C7436 XA1.XA4.MN0.G a_3440_41636# 6.69e-20
C7437 XA20.XA2.MN1.D a_22448_44100# 8.29e-20
C7438 a_4808_51140# a_4808_50788# 0.0109f
C7439 D<7> D<4> 0.00124f
C7440 a_17408_51140# D<1> 0.0688f
C7441 AVDD XA4.XA3.MN0.G 2.47f
C7442 XA1.XA7.MP0.D a_3440_50084# 7.44e-20
C7443 D<6> D<5> 0.832f
C7444 XA0.XA6.MP2.G D<3> 8.62e-19
C7445 XB2.XA4.MP0.D m3_16544_1364# 0.0634f
C7446 XB1.XA3.MN1.D m3_7544_308# 0.0137f
C7447 EN XA2.XA1.XA4.MN0.D 3.17e-19
C7448 XA4.XA1.XA5.MP0.D a_11000_43044# 0.00176f
C7449 XA8.XA1.XA5.MP0.D a_21080_43396# 0.049f
C7450 XA3.XA3.MN0.G a_8480_40228# 0.00307f
C7451 a_19928_50084# a_21080_50084# 0.00133f
C7452 a_7328_50084# a_7328_49732# 0.0109f
C7453 XA7.XA6.MP0.G VREF 0.568f
C7454 XA7.XA1.XA5.MN2.G a_16040_47972# 0.00363f
C7455 AVDD a_19928_43748# 0.00159f
C7456 XA6.XA6.MP0.G XA3.XA4.MN0.D 1.85e-19
C7457 D<8> li_14804_19596# 3.5e-20
C7458 SARP a_13808_2094# 2.97e-20
C7459 a_8480_42340# a_8480_41988# 0.0109f
C7460 XA3.XA1.XA5.MN2.G a_8480_44452# 5.11e-19
C7461 XA4.XA1.XA5.MN2.G a_7328_44452# 0.00486f
C7462 XA0.XA6.MP2.G a_920_44804# 2.36e-19
C7463 XA7.XA4.MN0.D a_18560_47268# 0.0963f
C7464 VREF a_2288_46916# 0.0536f
C7465 AVDD a_7328_41284# 0.361f
C7466 XA20.XA3a.MN0.G a_22448_46564# 0.0969f
C7467 a_13520_48324# a_14888_48324# 8.89e-19
C7468 a_2288_48324# XA1.XA4.MN0.G 0.0674f
C7469 AVDD a_2288_52900# 0.387f
C7470 XA2.XA12.MP0.G a_4808_53604# 0.1f
C7471 XA6.XA12.MP0.G XA7.XA12.MP0.G 0.00217f
C7472 XA3.XA11.MN1.G a_5960_53604# 0.0124f
C7473 XA7.XA11.MN1.G XA8.XA12.MP0.G 0.00122f
C7474 XA3.XA1.XA1.MP1.D a_7328_40580# 0.00176f
C7475 XA8.XA1.XA1.MN0.D a_19928_40932# 0.0535f
C7476 XA8.XA4.MN0.G XA7.XA1.XA5.MN2.D 0.0024f
C7477 XA7.XA4.MN0.G XA8.XA1.XA5.MN2.D 0.0024f
C7478 XA2.XA4.MN0.G a_4808_45156# 0.00865f
C7479 XA2.XA3.MN0.G a_4808_46564# 0.156f
C7480 a_16040_46916# a_16040_46564# 0.0109f
C7481 XA7.XA3.MN0.G XA8.XA3.MN0.G 0.0258f
C7482 XA7.XA1.XA5.MN2.G a_14888_42340# 3.12e-19
C7483 XA6.XA1.XA5.MN2.G a_16040_42340# 1.97e-19
C7484 XA4.XA10.MP0.G XA4.XA9.MN1.G 0.202f
C7485 XA20.XA10.MN1.D a_22448_51492# 1.97e-19
C7486 CK_SAMPLE XA2.XA6.MN2.D 0.0389f
C7487 AVDD a_14888_50788# 0.00154f
C7488 a_19928_52900# XA8.XA9.MN1.G 0.00113f
C7489 XB1.XA1.MP0.D a_8408_1742# 8.72e-20
C7490 a_13808_2446# XB2.XA4.MN0.D 0.00176f
C7491 a_14960_2446# XB2.M1.G 0.0696f
C7492 SAR_IP XB1.XA0.MP0.D 0.115f
C7493 XB1.M1.G XB1.XA4.MN0.D 0.139f
C7494 SAR_IN a_13808_2094# 0.00157f
C7495 a_9560_2446# a_9560_2094# 0.0109f
C7496 XA7.XA6.MP0.G XA7.XA1.XA1.MN0.D 0.00112f
C7497 SARN XDAC2.XC64b<1>.XRES1B.B 3.59f
C7498 XA20.XA3a.MN0.D XA0.XA1.XA4.MP1.D 0.0124f
C7499 a_4808_45156# a_4808_44804# 0.0109f
C7500 D<3> a_12368_39876# 7.77e-20
C7501 a_17408_45156# a_18560_45156# 0.00133f
C7502 XA4.XA4.MN0.G a_9848_42692# 0.0049f
C7503 XA1.XA3.MN0.G XA2.XA1.XA2.MP0.D 1.86e-19
C7504 a_12368_53252# VREF 0.00267f
C7505 AVDD a_17408_47972# 0.356f
C7506 XA0.XA9.MN1.G XA0.XA6.MP0.D 0.0618f
C7507 a_18560_51492# XA8.XA1.XA5.MN2.G 0.0658f
C7508 a_11000_51844# D<4> 1.25e-19
C7509 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES8.B 0.0228f
C7510 li_9184_26136# li_9184_25524# 0.00271f
C7511 XDAC1.XC64b<1>.XRES16.B XDAC1.X16ab.XRES16.B 0.0114f
C7512 XA20.XA2a.MN0.D XA3.XA1.XA1.MN0.S 0.137f
C7513 XA2.XA1.XA5.MP1.D a_5960_43396# 0.00176f
C7514 EN a_13520_43396# 0.00238f
C7515 AVDD a_4808_44452# 0.00125f
C7516 D<3> XA2.XA4.MN0.D 8.84e-19
C7517 D<2> XA0.XA4.MN0.D 0.0439f
C7518 a_7328_50436# a_7328_50084# 0.0109f
C7519 XDAC1.XC64a<0>.XRES2.B XDAC1.XC64a<0>.XRES16.B 0.457f
C7520 XDAC1.XC64a<0>.XRES8.B XDAC1.XC64a<0>.XRES1A.B 0.0228f
C7521 EN a_12368_40932# 0.00564f
C7522 XA0.XA1.XA4.MN0.D XA0.XA1.XA4.MP0.D 0.00918f
C7523 XA5.XA1.XA4.MP1.D a_12368_42340# 0.00176f
C7524 a_920_42692# a_920_42340# 0.0109f
C7525 D<0> a_21080_46564# 0.0695f
C7526 a_7328_49028# a_7328_48676# 0.0109f
C7527 XA0.XA6.MP2.G a_n232_45860# 0.0675f
C7528 XA4.XA1.XA5.MN2.G a_7328_45508# 0.00595f
C7529 XA3.XA1.XA5.MN2.G a_8480_45508# 9.01e-20
C7530 D<4> a_9848_46212# 0.0141f
C7531 D<1> XA20.XA2a.MN0.D 0.0858f
C7532 AVDD a_16040_42340# 0.361f
C7533 VREF XA1.XA4.MN0.G 0.263f
C7534 XA7.XA4.MN0.D a_17408_48324# 0.0682f
C7535 AVDD XA6.XA11.MN1.G 1.04f
C7536 a_23600_54308# CK_SAMPLE 0.0658f
C7537 a_11000_54308# a_11000_53956# 0.0109f
C7538 a_11000_41284# a_12368_41284# 8.89e-19
C7539 XA4.XA1.XA1.MN0.S XA4.XA1.XA1.MP1.D 0.0615f
C7540 SARP XDAC1.XC128a<1>.XRES1B.B 3.59f
C7541 XA2.XA1.XA5.MN2.G XA1.XA1.XA4.MN1.D 7.2e-19
C7542 XA20.XA10.MN1.D a_23600_40580# 0.0751f
C7543 D<1> XA7.XA1.XA2.MP0.D 0.0153f
C7544 a_2288_47268# a_2288_46916# 0.0109f
C7545 VREF a_3440_44804# 7.12e-19
C7546 XA1.XA4.MN0.D a_2288_44804# 9.15e-20
C7547 D<5> a_7328_43396# 7.77e-20
C7548 XA20.XA3a.MN0.D XA5.XA3.MN0.G 7.15e-20
C7549 XA5.XA4.MN0.G XA20.XA2a.MN0.D 0.00833f
C7550 XA1.XA4.MN0.G a_3440_46212# 0.0149f
C7551 XA8.XA4.MN0.G a_21080_46564# 3.46e-19
C7552 XA8.XA7.MP0.G a_19928_43044# 2.31e-19
C7553 XA0.XA12.MP0.D XA1.XA7.MP0.D 0.00283f
C7554 AVDD a_21080_51492# 0.387f
C7555 XA7.XA10.MP0.D a_17408_52900# 0.0877f
C7556 a_5960_52900# a_7328_52900# 8.89e-19
C7557 XA6.XA11.MN1.G a_13520_52196# 1.84e-19
C7558 a_21080_39876# a_22448_39876# 8.89e-19
C7559 XA20.XA3a.MN0.D a_21080_43748# 0.00346f
C7560 a_22448_45860# a_22448_45508# 0.0109f
C7561 XA6.XA4.MN0.G XA6.XA1.XA5.MP0.D 0.00138f
C7562 XA5.XA3.MN0.G a_12368_44452# 0.055f
C7563 XA8.XA1.XA5.MN2.G a_19928_40580# 0.083f
C7564 XA0.XA7.MP0.G a_3440_40228# 0.0825f
C7565 XA2.XA1.XA5.MN2.G a_2288_40228# 0.00255f
C7566 XA3.XA4.MN0.D XA3.XA1.XA4.MN0.D 8.11e-19
C7567 SARN a_12368_2094# 0.00496f
C7568 AVDD a_14888_49028# 0.00154f
C7569 a_5960_51844# XA2.XA8.MP0.D 0.0215f
C7570 a_16040_51844# a_17408_51844# 8.89e-19
C7571 CK_SAMPLE a_n232_49380# 0.00139f
C7572 D<5> li_9184_26136# 0.00504f
C7573 EN XA2.XA1.XA5.MP1.D 0.0544f
C7574 XA20.XA3a.MN0.D a_8480_41284# 0.00649f
C7575 XA20.XA2a.MN0.D XA7.XA1.XA4.MP0.D 0.0255f
C7576 XA1.XA3.MN0.G a_3440_41988# 0.00343f
C7577 XA3.XA8.MP0.D VREF 7.83e-19
C7578 D<4> XA2.XA6.MP0.G 0.0801f
C7579 D<3> XA1.XA6.MP0.G 0.11f
C7580 XA7.XA6.MN2.D a_18560_50436# 0.00176f
C7581 D<2> XA0.XA6.MP0.G 0.051f
C7582 AVDD a_4808_45508# 0.00131f
C7583 a_18560_50788# a_19928_50788# 8.89e-19
C7584 D<5> XA3.XA6.MP0.G 0.537f
C7585 a_4808_43044# a_4808_42692# 0.0109f
C7586 a_16040_43044# XA6.XA1.XA4.MP1.D 0.00176f
C7587 XA3.XA1.XA2.MP0.D a_8480_42340# 0.0966f
C7588 XA7.XA1.XA2.MP0.D XA7.XA1.XA4.MP0.D 4.34e-19
C7589 EN a_18560_41636# 1.25e-19
C7590 XA3.XA4.MN0.D a_8480_49380# 0.155f
C7591 VREF a_12368_49380# 0.0171f
C7592 AVDD a_23600_43044# 0.00181f
C7593 XA5.XA1.XA5.MN2.G XA4.XA3.MN0.G 0.106f
C7594 a_n232_49380# a_920_49380# 0.00133f
C7595 a_2288_41636# XA1.XA1.XA1.MN0.S 0.071f
C7596 D<2> a_14888_44100# 6.49e-19
C7597 a_8480_47972# a_8480_47620# 0.0109f
C7598 XA1.XA4.MN0.G a_2288_47268# 0.155f
C7599 XA0.XA7.MP0.G XA0.XA1.XA2.MP0.D 0.144f
C7600 XA7.XA4.MN0.D a_18560_46212# 1.1e-19
C7601 VREF a_2288_45860# 0.0178f
C7602 AVDD a_22448_40580# 0.483f
C7603 a_21080_47972# a_22448_47972# 8.89e-19
C7604 XA5.XA6.MP0.G a_12368_45156# 5.5e-19
C7605 XA20.XA12.MP0.G XA8.XA9.MN1.G 5.35e-19
C7606 XA3.XA11.MP0.D a_7328_53252# 0.0494f
C7607 XA5.XA11.MN1.G a_13520_52900# 0.00208f
C7608 a_8480_53604# XA3.XA10.MP0.D 1.17e-19
C7609 a_18560_53604# a_18560_53252# 0.0109f
C7610 AVDD a_3440_52196# 0.00154f
C7611 a_14888_40580# a_14888_40228# 0.0109f
C7612 XA4.XA1.XA5.MN2.G a_8480_41284# 0.00733f
C7613 VREF a_21080_43396# 3.39e-19
C7614 XA20.XA3.MN0.D a_23600_43044# 0.0828f
C7615 XA2.XA6.MP0.G XA2.XA1.XA4.MP0.D 9.97e-19
C7616 XA0.XA11.MN1.G a_12368_334# 0.00139f
C7617 a_14888_46212# a_16040_46212# 0.00133f
C7618 XA6.XA6.MP0.G a_16040_42692# 5.5e-19
C7619 XA5.XA3.MN0.G a_12368_45508# 0.0682f
C7620 XA8.XA9.MN0.D a_19928_52196# 0.0492f
C7621 XA8.XA9.MN1.G a_21080_52196# 0.0681f
C7622 AVDD a_14888_50084# 0.00144f
C7623 XA4.XA9.MN0.D XA4.XA7.MP0.D 0.00986f
C7624 CK_SAMPLE XA3.XA6.MP0.D 0.0278f
C7625 XA7.XA10.MP0.G XA7.XA8.MP0.D 0.0434f
C7626 XA2.XA10.MP0.G a_4808_51492# 6.8e-20
C7627 XA1.XA9.MN1.G a_2288_51844# 6.57e-19
C7628 a_12368_1038# a_12368_686# 0.0109f
C7629 XA6.XA6.MP0.G a_12368_39876# 0.00118f
C7630 a_8480_44452# a_9848_44452# 8.89e-19
C7631 XA2.XA1.XA5.MN2.D a_5960_43748# 0.00388f
C7632 XA8.XA1.XA5.MN2.D XA8.XA1.XA5.MP1.D 0.0488f
C7633 a_22448_44804# a_22448_44452# 0.0109f
C7634 a_21080_45156# EN 1.83e-19
C7635 SARN li_14804_19596# 0.00103f
C7636 XA6.XA1.XA5.MN2.G a_13520_50788# 1.87e-19
C7637 D<6> XA2.XA6.MP2.D 0.0399f
C7638 XA5.XA9.MN1.G a_13520_49732# 0.00119f
C7639 AVDD XA3.XA3.MN0.G 2.47f
C7640 XA0.XA9.MN1.G VREF 0.0732f
C7641 XB2.XA4.MP0.D m3_16472_1364# 0.106f
C7642 XB1.XA3.MN1.D m3_7472_308# 0.0137f
C7643 XDAC2.XC128b<2>.XRES2.B XDAC2.XC128b<2>.XRES16.B 0.457f
C7644 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128b<2>.XRES1A.B 0.0228f
C7645 XA0.XA6.MP0.G XDAC2.XC32a<0>.XRES2.B 2.23e-21
C7646 EN XA1.XA1.XA4.MN0.D 3.17e-19
C7647 XA20.XA2a.MN0.D a_n232_40580# 0.00139f
C7648 XA8.XA1.XA5.MP0.D a_19928_43396# 2.16e-19
C7649 XA8.XA1.XA5.MN0.D a_21080_43396# 2.16e-19
C7650 a_8480_43396# a_9848_43396# 8.89e-19
C7651 XA3.XA4.MN0.D li_9184_24912# 0.00504f
C7652 XA6.XA6.MP0.D VREF 0.0115f
C7653 XA2.XA6.MP0.G a_5960_49380# 0.0781f
C7654 XA5.XA6.MP0.G XA5.XA4.MN0.D 0.76f
C7655 XA8.XA6.MN0.D a_19928_49732# 0.00176f
C7656 XA8.XA6.MP0.G a_21080_49732# 0.101f
C7657 AVDD a_18560_43748# 0.00125f
C7658 SARP a_12368_2094# 0.0384f
C7659 a_19928_42340# a_21080_42340# 0.00133f
C7660 XA8.XA1.XA4.MN0.D a_19928_41988# 0.00176f
C7661 a_7328_42692# XA3.XA1.XA1.MN0.S 6.76e-20
C7662 XA8.XA1.XA2.MP0.D a_21080_40932# 4.25e-20
C7663 XA7.XA4.MN0.D a_17408_47268# 0.0576f
C7664 VREF a_920_46916# 0.0536f
C7665 AVDD a_5960_41284# 0.361f
C7666 a_18560_48676# XA7.XA4.MN0.G 1.34e-19
C7667 XA0.XA6.MP2.G a_n232_44804# 5.24e-19
C7668 D<4> a_11000_45156# 6.68e-19
C7669 XA3.XA1.XA5.MN2.G a_7328_44452# 7.1e-20
C7670 XA4.XA1.XA5.MN2.G a_5960_44452# 7.1e-20
C7671 CK_SAMPLE XA8.XA11.MP0.D 0.0011f
C7672 AVDD a_920_52900# 0.387f
C7673 a_17408_53956# a_17408_53604# 0.0109f
C7674 XA7.XA11.MN1.G XA7.XA12.MP0.G 0.278f
C7675 XA3.XA11.MN1.G a_4808_53604# 0.00305f
C7676 XA6.XA12.MP0.G XA8.XA11.MN1.G 1.54e-19
C7677 SARP li_9184_9156# 0.00103f
C7678 XA2.XA1.XA1.MN0.S a_5960_39876# 2.54e-19
C7679 XA7.XA1.XA1.MN0.S a_18560_40228# 0.0215f
C7680 a_7328_40932# a_8480_40932# 0.00133f
C7681 XA2.XA4.MN0.G a_3440_45156# 2.2e-19
C7682 XA1.XA4.MN0.G a_4808_45156# 2.2e-19
C7683 XA7.XA4.MN0.G XA7.XA1.XA5.MN2.D 0.135f
C7684 XA6.XA1.XA5.MN2.G a_14888_42340# 0.00568f
C7685 XA0.XA11.MN1.G a_13808_3854# 0.00283f
C7686 a_n232_52548# XA0.XA9.MN0.D 0.00176f
C7687 a_920_52548# XA0.XA9.MN1.G 0.0658f
C7688 a_12368_52548# a_13520_52548# 0.00133f
C7689 CK_SAMPLE D<6> 0.0523f
C7690 AVDD a_13520_50788# 0.00154f
C7691 XB2.XA1.MN0.D a_13808_2094# 4.63e-19
C7692 XB1.XA1.MN0.D XB1.XA0.MP0.D 0.0115f
C7693 a_13808_2446# XB2.M1.G 0.0339f
C7694 XB1.M1.G XB1.XA4.MP0.D 0.233f
C7695 SAR_IN a_12368_2094# 0.0503f
C7696 a_14960_3502# XB2.XA3.MN1.D 1.93e-19
C7697 XA20.XA3a.MN0.D XA0.XA1.XA4.MN1.D 0.0124f
C7698 XA5.XA1.XA5.MN2.D a_13520_44804# 0.153f
C7699 a_11000_53252# VREF 0.00292f
C7700 XA0.XA9.MN1.G XA0.XA6.MN0.D 0.0615f
C7701 AVDD a_16040_47972# 0.356f
C7702 a_7328_51492# a_7328_51140# 0.0109f
C7703 a_17408_51492# XA8.XA1.XA5.MN2.G 0.0714f
C7704 XA5.XA9.MN1.G a_13520_50436# 0.01f
C7705 XA0.XA7.MP0.G XA2.XA1.XA5.MN2.G 1.58f
C7706 a_8480_43748# XA3.XA1.XA5.MN0.D 0.00176f
C7707 XA7.XA1.XA5.MP1.D XA7.XA1.XA5.MP0.D 0.0488f
C7708 XA7.XA1.XA5.MN1.D XA7.XA1.XA2.MP0.D 0.0102f
C7709 XA20.XA2a.MN0.D XA2.XA1.XA1.MP2.D 0.0102f
C7710 EN a_12368_43396# 0.162f
C7711 AVDD a_3440_44452# 0.00125f
C7712 XA3.XA6.MP0.G XA4.XA6.MP0.G 4.3f
C7713 XA2.XA6.MP0.G XA5.XA6.MP0.G 0.0325f
C7714 a_21080_50436# XA8.XA6.MP0.G 0.0662f
C7715 a_19928_50436# XA8.XA6.MN0.D 0.00176f
C7716 XA5.XA6.MP2.D VREF 5.13e-19
C7717 D<3> XA1.XA4.MN0.D 0.0332f
C7718 D<4> XA4.XA4.MN0.D 0.203f
C7719 XA0.XA6.MP0.G XA7.XA6.MP0.G 0.0811f
C7720 XA1.XA6.MP0.G XA6.XA6.MP0.G 0.0781f
C7721 EN a_11000_40932# 0.00564f
C7722 a_12368_42692# XA5.XA1.XA4.MP0.D 0.00176f
C7723 D<8> li_14804_30036# 0.00508f
C7724 D<0> a_19928_46564# 0.0551f
C7725 a_18560_49028# a_19928_49028# 8.89e-19
C7726 XA3.XA1.XA5.MN2.G a_7328_45508# 7.1e-20
C7727 XA4.XA1.XA5.MN2.G a_5960_45508# 7.1e-20
C7728 XA20.XA10.MN1.D a_23600_43044# 0.00386f
C7729 AVDD a_14888_42340# 0.00125f
C7730 VREF XA0.XA4.MN0.G 0.263f
C7731 DONE a_23600_53956# 2.14e-19
C7732 XA20.XA11.MP0.D a_22448_53956# 0.00176f
C7733 a_22448_54308# CK_SAMPLE 0.0734f
C7734 AVDD XA4.XA12.MP0.G 0.709f
C7735 XA20.XA1.MN0.D a_23600_40228# 0.00339f
C7736 XA4.XA1.XA1.MN0.S XA4.XA1.XA1.MN0.D 0.0743f
C7737 XA2.XA1.XA5.MN2.G XA1.XA1.XA4.MP1.D 0.00353f
C7738 XA0.XA7.MP0.G XA1.XA1.XA4.MN1.D 0.0131f
C7739 XA20.XA10.MN1.D a_22448_40580# 0.0676f
C7740 VREF a_2288_44804# 0.0691f
C7741 XA20.XA3a.MN0.D XA4.XA3.MN0.G 7.15e-20
C7742 XA4.XA4.MN0.G XA20.XA2a.MN0.D 0.00823f
C7743 XA8.XA4.MN0.G a_19928_46564# 0.0155f
C7744 XA1.XA4.MN0.G a_2288_46212# 3.46e-19
C7745 a_13520_47268# a_14888_47268# 8.89e-19
C7746 XA8.XA1.XA5.MN2.G a_19928_43044# 0.0748f
C7747 AVDD a_19928_51492# 0.00166f
C7748 XA0.XA11.MN1.G XA0.XA9.MN1.G 0.00804f
C7749 XA0.XA12.MP0.D XA0.XA7.MP0.D 8.25e-19
C7750 CK_SAMPLE a_14888_51844# 1.64e-19
C7751 XA0.XA10.MP0.D XA0.XA10.MP0.G 0.194f
C7752 XA20.XA3a.MN0.D a_19928_43748# 0.00352f
C7753 XA6.XA4.MN0.G XA6.XA1.XA5.MN0.D 0.0198f
C7754 a_8480_45508# a_9848_45508# 8.89e-19
C7755 a_12368_45860# XA5.XA1.XA5.MN2.D 3.12e-20
C7756 XA7.XA1.XA5.MN2.G a_19928_40580# 7.1e-20
C7757 XA8.XA1.XA5.MN2.G a_18560_40580# 0.00564f
C7758 XA0.XA7.MP0.G a_2288_40228# 0.0128f
C7759 XA3.XA4.MN0.D XA3.XA1.XA4.MP0.D 7.97e-19
C7760 SARN a_11000_2094# 0.0413f
C7761 XA4.XA9.MN1.G a_11000_51140# 0.0222f
C7762 AVDD a_13520_49028# 0.00154f
C7763 a_4808_51844# XA2.XA8.MP0.D 0.0215f
C7764 XA2.XA7.MP0.D a_5960_51492# 0.0893f
C7765 CK_SAMPLE XA8.XA4.MN0.D 0.027f
C7766 a_5960_52196# XA3.XA1.XA5.MN2.G 3.39e-19
C7767 XDAC1.XC0.XRES4.B XDAC1.XC64b<1>.XRES4.B 0.00284f
C7768 li_9184_31260# li_9184_30648# 0.00271f
C7769 XDAC1.XC0.XRES2.B XDAC1.XC0.XRES1A.B 0.0136f
C7770 a_3440_44100# a_3440_43748# 0.0109f
C7771 a_14888_44100# XA6.XA1.XA5.MN1.D 0.00176f
C7772 EN XA2.XA1.XA5.MN1.D 0.0157f
C7773 XA20.XA2a.MN0.D XA6.XA1.XA4.MP0.D 0.0251f
C7774 XA3.XA1.XA5.MN2.D a_8480_43044# 5.1e-20
C7775 a_3440_44452# XA1.XA1.XA2.MP0.D 5.16e-20
C7776 XA0.XA6.MP2.G li_9184_24912# 3.5e-20
C7777 SARN XDAC2.XC64a<0>.XRES1A.B 3.59f
C7778 XA2.XA8.MP0.D VREF 7.83e-19
C7779 a_5960_50788# a_5960_50436# 0.0109f
C7780 AVDD a_3440_45508# 0.00131f
C7781 XDAC1.XC32a<0>.XRES1B.B XDAC1.XC32a<0>.XRES4.B 0.428f
C7782 XA1.XA1.XA4.MP1.D XA1.XA1.XA4.MN1.D 0.00918f
C7783 XA3.XA1.XA2.MP0.D a_7328_42340# 2.54e-19
C7784 XA0.XA4.MN0.D XDAC1.XC32a<0>.XRES2.B 2.23e-21
C7785 EN a_17408_41636# 0.00649f
C7786 a_18560_49732# a_18560_49380# 0.0109f
C7787 XA3.XA4.MN0.D a_7328_49380# 0.154f
C7788 VREF a_11000_49380# 0.0171f
C7789 XA4.XA6.MP0.G a_11000_48324# 0.00417f
C7790 AVDD a_22448_43044# 0.419f
C7791 XA5.XA1.XA5.MN2.G XA3.XA3.MN0.G 0.0021f
C7792 XA4.XA1.XA5.MN2.G XA4.XA3.MN0.G 5.78e-19
C7793 XA8.XA6.MP0.G a_21080_48676# 0.0881f
C7794 a_13520_41636# a_14888_41636# 8.89e-19
C7795 SARP XDAC1.XC64b<1>.XRES1B.B 3.59f
C7796 D<5> EN 0.0614f
C7797 XA7.XA4.MN0.G a_18560_47620# 0.154f
C7798 XA7.XA1.XA5.MN2.G a_16040_43748# 0.00442f
C7799 VREF a_920_45860# 0.0178f
C7800 AVDD a_21080_40580# 0.381f
C7801 XA4.XA12.MP0.G a_11000_52900# 1.28e-19
C7802 XA5.XA11.MN1.G a_12368_52900# 0.00273f
C7803 AVDD a_2288_52196# 0.37f
C7804 a_920_40228# a_2288_40228# 8.89e-19
C7805 XA4.XA4.MN0.G a_11000_44100# 6.11e-19
C7806 XA20.XA3.MN0.D a_22448_43044# 0.00246f
C7807 XA2.XA6.MP0.G XA2.XA1.XA4.MN0.D 6.07e-19
C7808 XA0.XA11.MN1.G a_11000_334# 0.00139f
C7809 a_2288_46212# a_2288_45860# 0.0109f
C7810 XA6.XA6.MP0.G a_14888_42692# 7.76e-20
C7811 XA3.XA1.XA5.MN2.G a_8480_41284# 0.00392f
C7812 XA4.XA1.XA5.MN2.G a_7328_41284# 0.0169f
C7813 XA8.XA9.MN1.G a_19928_52196# 0.0862f
C7814 AVDD a_13520_50084# 0.00144f
C7815 XA4.XA9.MN1.G XA4.XA7.MP0.D 0.274f
C7816 a_7328_52196# a_8480_52196# 0.00133f
C7817 CK_SAMPLE XA3.XA6.MP0.G 0.0463f
C7818 XB2.XA3.MN1.D a_14960_334# 0.00886f
C7819 XB1.XA3.MN1.D a_9560_n18# 9.07e-19
C7820 XA7.XA4.MN0.G a_18560_41988# 1.74e-19
C7821 XA20.XA2a.MN0.D a_n232_43044# 1.43e-19
C7822 XA2.XA1.XA5.MN2.D a_4808_43748# 0.00224f
C7823 XA8.XA1.XA5.MN2.D XA8.XA1.XA5.MN1.D 0.0488f
C7824 a_19928_45156# EN 4.58e-19
C7825 XA6.XA1.XA5.MN2.G a_12368_50788# 0.00548f
C7826 a_3440_51140# a_3440_50788# 0.0109f
C7827 D<6> XA2.XA6.MN2.D 1.59e-19
C7828 XA5.XA9.MN1.G a_12368_49732# 0.0215f
C7829 AVDD XA2.XA3.MN0.G 2.47f
C7830 XA0.XA9.MN1.G XA0.XA4.MN0.D 0.00938f
C7831 a_16040_51140# XA6.XA6.MP2.D 0.00176f
C7832 XB2.XA4.MP0.D m3_26048_2244# 0.0273f
C7833 XB1.XA3.MN1.D m3_n1960_1188# 0.0634f
C7834 EN XA1.XA1.XA4.MP0.D 0.0386f
C7835 XA4.XA1.XA2.MP0.D a_11000_43044# 3.59e-19
C7836 XA0.XA1.XA2.MP0.D XA0.XA1.XA4.MP1.D 4.34e-19
C7837 XA4.XA1.XA5.MN0.D a_9848_43044# 0.00176f
C7838 XA8.XA1.XA5.MN0.D a_19928_43396# 0.0474f
C7839 a_18560_50084# a_19928_50084# 8.89e-19
C7840 a_5960_50084# a_5960_49732# 0.0109f
C7841 XA2.XA6.MP0.G a_4808_49380# 0.0547f
C7842 XA8.XA6.MP0.G a_19928_49732# 0.00239f
C7843 AVDD a_17408_43748# 0.357f
C7844 D<8> XDAC2.XC128b<2>.XRES1A.B 4.06e-21
C7845 SARP a_11000_2094# 0.00802f
C7846 a_7328_42340# a_7328_41988# 0.0109f
C7847 XA0.XA4.MN0.D a_920_46916# 0.00254f
C7848 AVDD a_4808_41284# 0.00125f
C7849 a_12368_48324# a_13520_48324# 0.00133f
C7850 a_920_48324# XA0.XA4.MN0.G 0.0658f
C7851 D<4> a_9848_45156# 7.77e-19
C7852 XA3.XA1.XA5.MN2.G a_5960_44452# 0.00486f
C7853 AVDD a_n232_52900# 0.00166f
C7854 XA7.XA11.MN1.G XA8.XA11.MN1.G 0.271f
C7855 XA2.XA11.MN1.G a_5960_53604# 0.0658f
C7856 XA2.XA1.XA1.MN0.S a_4808_39876# 2.54e-19
C7857 XA7.XA1.XA1.MN0.S a_17408_40228# 0.0313f
C7858 XA2.XA1.XA1.MP1.D a_5960_40580# 0.00176f
C7859 XA7.XA1.XA1.MN0.D a_18560_40932# 0.0535f
C7860 a_14888_46916# a_14888_46564# 0.0109f
C7861 XA1.XA3.MN0.G a_3440_46564# 0.156f
C7862 XA1.XA4.MN0.G a_3440_45156# 0.00865f
C7863 D<3> a_13520_42692# 6.49e-19
C7864 XA6.XA3.MN0.G XA7.XA3.MN0.G 0.00869f
C7865 D<7> XA1.XA1.XA4.MN0.D 0.00144f
C7866 XA6.XA1.XA5.MN2.G a_13520_42340# 4.69e-19
C7867 XA7.XA6.MP0.G XA7.XA1.XA5.MN0.D 7.41e-19
C7868 XA3.XA4.MN0.D XA3.XA1.XA5.MN1.D 9.89e-19
C7869 VREF XA5.XA1.XA5.MP1.D 0.00623f
C7870 XA0.XA11.MN1.G a_9560_3150# 0.0101f
C7871 a_n232_52548# XA0.XA9.MN1.G 0.0727f
C7872 CK_SAMPLE XA1.XA6.MN2.D 0.0389f
C7873 AVDD a_12368_50788# 0.363f
C7874 XA3.XA10.MP0.G XA3.XA9.MN0.D 0.106f
C7875 a_12368_2446# XB2.M1.G 1.17e-19
C7876 XB1.XA1.MP0.D XB1.XA0.MP0.D 0.0524f
C7877 a_8408_2446# a_8408_2094# 0.0109f
C7878 SARN li_14804_30036# 0.00103f
C7879 XA5.XA1.XA5.MN2.D a_12368_44804# 0.156f
C7880 a_3440_45156# a_3440_44804# 0.0109f
C7881 a_16040_45156# a_17408_45156# 8.89e-19
C7882 XA3.XA6.MP0.G a_8480_40932# 3.97e-20
C7883 XA3.XA4.MN0.G a_8480_42692# 0.0049f
C7884 XA2.XA3.MN0.G XA1.XA1.XA2.MP0.D 0.00181f
C7885 XA0.XA9.MN1.G XA0.XA6.MP0.G 0.0725f
C7886 AVDD a_14888_47972# 0.00125f
C7887 XA5.XA9.MN1.G a_12368_50436# 7.76e-19
C7888 XA7.XA7.MP0.D D<1> 2.65e-19
C7889 XDAC2.X16ab.XRES1B.B XDAC2.X16ab.XRES4.B 0.428f
C7890 a_22448_43748# a_23600_43748# 0.00133f
C7891 XA7.XA1.XA5.MP1.D XA7.XA1.XA2.MP0.D 6.52e-20
C7892 XA20.XA2a.MN0.D XA2.XA1.XA1.MN0.S 0.137f
C7893 XA2.XA1.XA5.MN1.D a_4808_43396# 0.00176f
C7894 EN a_11000_43396# 0.162f
C7895 a_19928_50436# XA8.XA6.MP0.G 3.02e-20
C7896 D<3> VREF 1.3f
C7897 XA6.XA1.XA5.MN2.G a_12368_49028# 0.00363f
C7898 AVDD a_2288_44452# 0.357f
C7899 D<7> a_3440_49380# 5.91e-19
C7900 D<4> XA3.XA4.MN0.D 3.22f
C7901 D<1> a_18560_49732# 7.01e-19
C7902 a_5960_50436# a_5960_50084# 0.0109f
C7903 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC1.XRES1B.B 0.00444f
C7904 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES1A.B 0.0197f
C7905 li_14804_10992# li_14804_10380# 0.00271f
C7906 XDAC2.XC64a<0>.XRES8.B XDAC2.XC64a<0>.XRES16.B 0.0904f
C7907 XA5.XA1.XA2.MP0.D XA5.XA1.XA1.MN0.S 2.11e-19
C7908 XA4.XA1.XA4.MP1.D a_11000_42340# 0.00176f
C7909 a_n232_42692# a_n232_42340# 0.0109f
C7910 XA8.XA6.MP0.G a_21080_47620# 8.5e-20
C7911 a_5960_49028# a_5960_48676# 0.0109f
C7912 XA3.XA1.XA5.MN2.G a_5960_45508# 0.00595f
C7913 AVDD a_13520_42340# 0.00125f
C7914 XA4.XA6.MP0.G a_11000_47268# 5.95e-19
C7915 XA6.XA4.MN0.D a_16040_48324# 0.0698f
C7916 XA0.XA4.MN0.D XA0.XA4.MN0.G 0.728f
C7917 XA0.XA6.MP0.G a_920_46916# 5.5e-19
C7918 XA20.XA11.MN0.D a_23600_53956# 0.0316f
C7919 DONE a_22448_53956# 0.00574f
C7920 a_9848_54308# a_9848_53956# 0.0109f
C7921 a_22448_54308# a_23600_54308# 0.00133f
C7922 AVDD XA5.XA11.MN1.G 1.89f
C7923 a_9848_41284# a_11000_41284# 0.00133f
C7924 XA20.XA1.MN0.D a_22448_40228# 0.0215f
C7925 SARP li_9184_19596# 0.00103f
C7926 VREF a_920_44804# 0.0691f
C7927 XA0.XA7.MP0.G XA1.XA1.XA4.MP1.D 7.44e-19
C7928 XA4.XA6.MP0.G EN 0.071f
C7929 XA20.XA3a.MN0.D XA3.XA3.MN0.G 0.223f
C7930 XA2.XA6.MP0.G XA2.XA1.XA5.MP1.D 0.00121f
C7931 XA3.XA4.MN0.G XA20.XA2a.MN0.D 0.00833f
C7932 XA7.XA4.MN0.G a_19928_46564# 2.2e-19
C7933 XA8.XA4.MN0.G a_18560_46564# 2.2e-19
C7934 AVDD a_9560_2446# 0.00166f
C7935 a_920_47268# a_920_46916# 0.0109f
C7936 XA8.XA1.XA5.MN2.G a_18560_43044# 2.31e-19
C7937 CK_SAMPLE a_13520_51844# 2.08e-19
C7938 AVDD a_18560_51492# 0.00166f
C7939 XA5.XA11.MN1.G a_13520_52196# 5.56e-19
C7940 XA6.XA10.MP0.D a_16040_52900# 0.0893f
C7941 a_4808_52900# a_5960_52900# 0.00133f
C7942 a_19928_39876# a_21080_39876# 0.00133f
C7943 XA4.XA3.MN0.G a_11000_44452# 0.055f
C7944 XA6.XA4.MN0.G XA6.XA1.XA2.MP0.D 0.206f
C7945 a_21080_45860# a_21080_45508# 0.0109f
C7946 XA7.XA1.XA5.MN2.G a_18560_40580# 0.0806f
C7947 XA8.XA1.XA5.MN2.G a_17408_40580# 0.0431f
C7948 XA0.XA7.MP0.G a_920_40228# 0.0108f
C7949 XA4.XA6.MP0.G a_11000_41636# 5.5e-19
C7950 D<2> XA6.XA1.XA1.MN0.D 0.0192f
C7951 SARN a_9560_2094# 2.97e-20
C7952 XA20.XA3a.MN0.D a_18560_43748# 0.00228f
C7953 XA4.XA9.MN1.G a_9848_51140# 0.0469f
C7954 AVDD a_12368_49028# 0.356f
C7955 XA7.XA7.MP0.D XA7.XA8.MP0.D 0.124f
C7956 a_14888_51844# a_16040_51844# 0.00133f
C7957 XA2.XA7.MP0.D a_4808_51492# 0.124f
C7958 CK_SAMPLE XA7.XA4.MN0.D 0.0364f
C7959 a_7328_53956# VREF 0.00396f
C7960 D<5> XDAC1.X16ab.XRES1B.B 0.00405f
C7961 EN XA1.XA1.XA5.MN1.D 0.0157f
C7962 XA20.XA2a.MN0.D XA6.XA1.XA4.MN0.D 0.0375f
C7963 XA3.XA1.XA5.MN2.D a_7328_43044# 1.88e-19
C7964 a_13520_44804# XA5.XA1.XA2.MP0.D 2.6e-20
C7965 XA1.XA8.MP0.D VREF 7.83e-19
C7966 D<1> a_18560_50436# 5.7e-19
C7967 XA7.XA6.MP2.D a_17408_50436# 0.00176f
C7968 AVDD a_2288_45508# 0.359f
C7969 a_17408_50788# a_18560_50788# 0.00133f
C7970 XA6.XA1.XA5.MN2.G a_12368_50084# 0.00366f
C7971 a_3440_43044# a_3440_42692# 0.0109f
C7972 a_14888_43044# XA6.XA1.XA4.MN1.D 0.00176f
C7973 EN a_16040_41636# 0.00649f
C7974 XA4.XA1.XA5.MN2.G XA3.XA3.MN0.G 0.225f
C7975 XA8.XA7.MP0.G a_22448_46916# 6.64e-19
C7976 VREF a_9848_49380# 8.08e-19
C7977 XA4.XA6.MP0.G a_9848_48324# 0.00295f
C7978 AVDD a_21080_43044# 0.381f
C7979 XA0.XA6.MP0.G XA0.XA4.MN0.G 0.0408f
C7980 XA8.XA6.MP0.G a_19928_48676# 0.0651f
C7981 a_920_41636# XA0.XA1.XA1.MP2.D 0.00176f
C7982 a_7328_47972# a_7328_47620# 0.0109f
C7983 XA0.XA4.MN0.G a_920_47268# 0.155f
C7984 XA7.XA4.MN0.G a_17408_47620# 0.155f
C7985 XA7.XA1.XA5.MN2.G a_14888_43748# 1.95e-19
C7986 XA0.XA4.MN0.D a_920_45860# 9.14e-20
C7987 VREF a_n232_45860# 1.19e-19
C7988 AVDD a_19928_40580# 0.00154f
C7989 a_19928_47972# a_21080_47972# 0.00133f
C7990 XA2.XA11.MP0.D a_5960_53252# 0.0494f
C7991 XA4.XA12.MP0.G a_9848_52900# 0.00258f
C7992 XA5.XA11.MN1.G a_11000_52900# 0.00183f
C7993 a_17408_53604# a_17408_53252# 0.0109f
C7994 AVDD a_920_52196# 0.37f
C7995 a_13520_40580# a_13520_40228# 0.0109f
C7996 XA4.XA4.MN0.G a_9848_44100# 0.0164f
C7997 XA0.XA11.MN1.G a_9560_334# 0.00214f
C7998 XA20.XA3a.MN0.D a_3440_44452# 2.59e-20
C7999 a_13520_46212# a_14888_46212# 8.89e-19
C8000 XA4.XA3.MN0.G a_11000_45508# 0.0698f
C8001 XA3.XA1.XA5.MN2.G a_7328_41284# 5.96e-19
C8002 XA8.XA9.MN1.G a_18560_52196# 2.84e-19
C8003 AVDD a_12368_50084# 0.358f
C8004 XA4.XA9.MN1.G XA3.XA7.MP0.D 0.00108f
C8005 CK_SAMPLE XA2.XA6.MP0.D 0.0276f
C8006 XA6.XA10.MP0.G XA6.XA8.MP0.D 0.0434f
C8007 XA1.XA10.MP0.G a_3440_51492# 6.8e-20
C8008 a_13808_1390# CK_SAMPLE_BSSW 2.9e-19
C8009 a_11000_1038# a_11000_686# 0.0109f
C8010 XB1.XA3.MN1.D a_8408_n18# 0.0124f
C8011 XB2.XA3.MN1.D a_13808_334# 9.07e-19
C8012 XA7.XA4.MN0.G a_17408_41988# 5.1e-20
C8013 a_7328_44452# a_8480_44452# 0.00133f
C8014 XA20.XA2a.MN0.D a_23600_43396# 0.00246f
C8015 a_21080_44804# a_21080_44452# 0.0109f
C8016 a_18560_45156# EN 4.58e-19
C8017 SARN XDAC2.XC128b<2>.XRES1A.B 3.59f
C8018 XA5.XA6.MP0.G a_13520_39876# 7.76e-20
C8019 XA20.XA3a.MN0.D a_14888_42340# 0.00547f
C8020 AVDD XA1.XA3.MN0.G 2.47f
C8021 XA5.XA1.XA5.MN2.G a_12368_50788# 7.1e-20
C8022 XA6.XA1.XA5.MN2.G a_11000_50788# 7.1e-20
C8023 XA0.XA6.MP2.G D<4> 0.0013f
C8024 a_22448_52548# VREF 0.00104f
C8025 D<7> D<5> 0.146f
C8026 XB1.XA3.MN1.D m3_n2104_1188# 0.17f
C8027 XB2.XA4.MP0.D m3_25976_2244# 0.0137f
C8028 XDAC1.XC128b<2>.XRES2.B XDAC1.XC128b<2>.XRES16.B 0.457f
C8029 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128b<2>.XRES1A.B 0.0228f
C8030 XA0.XA6.MP0.G li_14804_14472# 1.85e-20
C8031 XA20.XA2a.MN0.D a_22448_40932# 6.25e-19
C8032 XA0.XA1.XA2.MP0.D XA0.XA1.XA4.MN1.D 0.056f
C8033 XA4.XA1.XA2.MP0.D a_9848_43044# 0.0292f
C8034 a_7328_43396# a_8480_43396# 0.00133f
C8035 XA8.XA1.XA2.MP0.D a_19928_43396# 0.0945f
C8036 XA3.XA4.MN0.D XDAC1.X16ab.XRES8.B 0.00669f
C8037 EN XA0.XA1.XA4.MP0.D 0.0392f
C8038 D<1> a_18560_48676# 3.48e-19
C8039 AVDD a_16040_43748# 0.357f
C8040 XA6.XA6.MP0.G VREF 0.568f
C8041 D<5> a_8480_48324# 6.53e-19
C8042 SARP a_9560_2094# 0.00112f
C8043 a_18560_42340# a_19928_42340# 8.89e-19
C8044 XA7.XA1.XA4.MN0.D a_18560_41988# 0.00176f
C8045 XA4.XA6.MP0.G a_11000_46212# 5.5e-19
C8046 XA0.XA6.MP0.G a_920_45860# 5.5e-19
C8047 XA6.XA4.MN0.D a_16040_47268# 0.0576f
C8048 XA0.XA4.MN0.D a_n232_46916# 0.00456f
C8049 AVDD a_3440_41284# 0.00125f
C8050 a_n232_48324# XA0.XA4.MN0.G 0.0677f
C8051 XA3.XA1.XA5.MN2.G a_4808_44452# 1.86e-19
C8052 D<1> XA7.XA1.XA5.MN2.D 0.0348f
C8053 AVDD XA20.XA9.MP0.D 4.02f
C8054 XA7.XA11.MN1.G XA6.XA12.MP0.G 0.142f
C8055 DONE a_23600_53252# 2.31e-19
C8056 a_16040_53956# a_16040_53604# 0.0109f
C8057 XA1.XA12.MP0.G a_3440_53604# 0.102f
C8058 XA2.XA11.MN1.G a_4808_53604# 0.0709f
C8059 SARP XDAC1.XC64a<0>.XRES1A.B 3.59f
C8060 XA2.XA1.XA1.MN0.D a_5960_40580# 8.3e-19
C8061 XA7.XA1.XA1.MN0.D a_17408_40932# 8.29e-20
C8062 a_5960_40932# a_7328_40932# 8.89e-19
C8063 XA1.XA3.MN0.G a_2288_46564# 0.155f
C8064 XA1.XA4.MN0.G a_2288_45156# 5.54e-19
C8065 XA6.XA4.MN0.G XA6.XA1.XA5.MN2.D 0.135f
C8066 XA3.XA6.MP0.G a_8480_43396# 7.76e-20
C8067 D<3> a_12368_42692# 7.77e-20
C8068 D<7> XA1.XA1.XA4.MP0.D 6.09e-19
C8069 XA5.XA1.XA5.MN2.G a_13520_42340# 0.00568f
C8070 XA6.XA1.XA5.MN2.G a_12368_42340# 0.00442f
C8071 XA7.XA6.MP0.G XA7.XA1.XA5.MP0.D 0.00121f
C8072 XA3.XA4.MN0.D XA3.XA1.XA5.MP1.D 9.71e-19
C8073 VREF XA4.XA1.XA5.MP1.D 0.00623f
C8074 a_11000_52548# a_12368_52548# 8.89e-19
C8075 a_18560_52900# XA7.XA9.MN1.G 0.00113f
C8076 CK_SAMPLE XA1.XA6.MP2.D 3.06e-19
C8077 AVDD a_11000_50788# 0.363f
C8078 XA3.XA10.MP0.G XA3.XA9.MN1.G 0.202f
C8079 DONE XA8.XA6.MP2.D 2.25e-19
C8080 a_14960_3854# XB2.XA3.MN1.D 1.93e-19
C8081 XA0.XA4.MN0.D XA0.XA1.XA1.MN0.S 0.0163f
C8082 XA7.XA6.MP0.G XA6.XA1.XA1.MN0.D 4.63e-19
C8083 XA20.XA3a.MN0.D a_22448_43044# 0.00246f
C8084 XA3.XA6.MP0.G a_7328_40932# 4.24e-19
C8085 XA3.XA4.MN0.G a_7328_42692# 0.00224f
C8086 XA8.XA3.MN0.G a_19928_43748# 2.78e-19
C8087 XA1.XA3.MN0.G XA1.XA1.XA2.MP0.D 0.0363f
C8088 AVDD a_13520_47972# 0.00125f
C8089 a_5960_51492# a_5960_51140# 0.0109f
C8090 a_16040_51492# XA7.XA1.XA5.MN2.G 0.0699f
C8091 XA0.XA7.MP0.D a_n232_50788# 3.29e-19
C8092 XA20.XA9.MP0.D XA20.XA3.MN0.D 0.35f
C8093 a_7328_43748# XA3.XA1.XA5.MP0.D 0.00176f
C8094 a_8480_43748# XA3.XA1.XA2.MP0.D 0.0686f
C8095 XA20.XA2a.MN0.D XA1.XA1.XA1.MP2.D 0.0102f
C8096 EN a_9848_43396# 0.00238f
C8097 XA20.XA3a.MN0.D a_21080_40580# 0.0674f
C8098 D<3> XA0.XA4.MN0.D 0.0441f
C8099 XA6.XA1.XA5.MN2.G a_11000_49028# 7.1e-20
C8100 XA5.XA1.XA5.MN2.G a_12368_49028# 7.1e-20
C8101 AVDD a_920_44452# 0.357f
C8102 D<7> a_2288_49380# 0.00891f
C8103 D<4> XA2.XA4.MN0.D 0.192f
C8104 XA4.XA6.MP2.D VREF 5.13e-19
C8105 D<1> a_17408_49732# 0.0109f
C8106 XA3.XA6.MP0.G XA3.XA6.MP0.D 0.0392f
C8107 a_11000_42692# XA4.XA1.XA4.MP0.D 0.00176f
C8108 D<8> XDAC2.XC0.XRES1A.B 0.00406f
C8109 a_17408_49028# a_18560_49028# 0.00133f
C8110 XA8.XA7.MP0.G a_22448_45860# 6.64e-19
C8111 XA3.XA1.XA5.MN2.G a_4808_45508# 2.31e-19
C8112 AVDD a_12368_42340# 0.361f
C8113 XA4.XA6.MP0.G a_9848_47268# 1.38e-19
C8114 VREF a_22448_48324# 0.00125f
C8115 XA6.XA4.MN0.D a_14888_48324# 0.0981f
C8116 D<2> XA20.XA2a.MN0.D 0.0851f
C8117 XA0.XA6.MP0.G a_n232_46916# 7.76e-20
C8118 DONE a_21080_53956# 0.00122f
C8119 XA20.XA11.MN0.D a_22448_53956# 3.74e-19
C8120 AVDD XA3.XA12.MP0.G 0.706f
C8121 XA8.XA1.XA1.MP2.D a_21080_41284# 0.0465f
C8122 VREF a_n232_44804# 7.12e-19
C8123 XA0.XA4.MN0.D a_920_44804# 9.14e-20
C8124 XA6.XA6.MP0.G a_16040_44100# 5.5e-19
C8125 XA0.XA7.MP0.G XA0.XA1.XA4.MP1.D 0.00353f
C8126 XA20.XA3a.MN0.D XA2.XA3.MN0.G 0.221f
C8127 XA2.XA6.MP0.G XA2.XA1.XA5.MN1.D 7.41e-19
C8128 XA2.XA4.MN0.G XA20.XA2a.MN0.D 0.00823f
C8129 XA7.XA4.MN0.G a_18560_46564# 0.0155f
C8130 XA0.XA4.MN0.G a_920_46212# 3.46e-19
C8131 AVDD a_8408_2446# 0.406f
C8132 a_12368_47268# a_13520_47268# 0.00133f
C8133 XA7.XA1.XA5.MN2.G a_18560_43044# 0.0732f
C8134 XA8.XA1.XA5.MN2.G a_17408_43044# 0.00551f
C8135 AVDD a_17408_51492# 0.387f
C8136 XA5.XA11.MN1.G a_12368_52196# 7.34e-19
C8137 a_23600_53252# a_23600_52900# 0.0109f
C8138 XA6.XA10.MP0.D a_14888_52900# 0.128f
C8139 a_7328_45508# a_8480_45508# 0.00133f
C8140 a_11000_45860# XA4.XA1.XA5.MN2.D 3.12e-20
C8141 XA4.XA3.MN0.G a_9848_44452# 0.0934f
C8142 D<6> a_5960_40932# 4.07e-20
C8143 XA7.XA1.XA5.MN2.G a_17408_40580# 0.00417f
C8144 XA0.XA7.MP0.G a_n232_40228# 5.59e-19
C8145 XA4.XA6.MP0.G a_9848_41636# 7.76e-20
C8146 XA2.XA4.MN0.D XA2.XA1.XA4.MP0.D 7.95e-19
C8147 XA0.XA6.MP0.G XA0.XA1.XA1.MN0.S 0.0143f
C8148 XA20.XA3a.MN0.D a_17408_43748# 0.00106f
C8149 AVDD a_11000_49028# 0.356f
C8150 XA20.XA9.MP0.D a_23600_50788# 0.00614f
C8151 a_3440_51844# XA1.XA8.MP0.D 0.0215f
C8152 CK_SAMPLE XA6.XA4.MN0.D 0.0364f
C8153 a_5960_53956# VREF 0.00366f
C8154 XA8.XA9.MN1.G XA8.XA7.MP0.G 0.049f
C8155 XA4.XA9.MN1.G a_8480_51140# 2.84e-19
C8156 XDAC2.XC0.XRES8.B XDAC2.XC0.XRES1A.B 0.0228f
C8157 XDAC2.XC0.XRES2.B XDAC2.XC0.XRES16.B 0.457f
C8158 XA0.XA1.XA5.MN1.D XA0.XA1.XA5.MP1.D 0.00918f
C8159 EN XA1.XA1.XA5.MP1.D 0.0543f
C8160 XA20.XA3a.MN0.D a_4808_41284# 0.00649f
C8161 XA20.XA2a.MN0.D XA5.XA1.XA4.MN0.D 0.0409f
C8162 XA0.XA6.MP2.G XDAC1.X16ab.XRES8.B 4.06e-21
C8163 SARN li_14804_9768# 0.00103f
C8164 a_13520_44100# XA5.XA1.XA5.MN1.D 0.00176f
C8165 a_2288_44100# a_2288_43748# 0.0109f
C8166 D<1> a_17408_50436# 0.0863f
C8167 a_4808_50788# a_4808_50436# 0.0109f
C8168 D<5> XA2.XA6.MP0.G 0.0629f
C8169 D<4> XA1.XA6.MP0.G 0.0801f
C8170 AVDD a_920_45508# 0.359f
C8171 D<3> XA0.XA6.MP0.G 0.102f
C8172 a_17408_51140# XA7.XA6.MP0.G 6.76e-20
C8173 XA6.XA1.XA5.MN2.G a_11000_50084# 7.1e-20
C8174 XA5.XA1.XA5.MN2.G a_12368_50084# 7.1e-20
C8175 XA0.XA8.MP0.D VREF 7.83e-19
C8176 XDAC2.XC128a<1>.XRES2.B XDAC2.XC32a<0>.XRES2.B 1.67e-19
C8177 li_14804_16116# li_14804_15696# 0.00411f
C8178 XA0.XA4.MN0.D li_9184_14472# 1.85e-20
C8179 EN a_14888_41636# 1.25e-19
C8180 XA4.XA1.XA5.MN2.G XA2.XA3.MN0.G 6.95e-19
C8181 XA3.XA1.XA5.MN2.G XA3.XA3.MN0.G 0.229f
C8182 XA8.XA7.MP0.G a_21080_46916# 0.00455f
C8183 VREF a_8480_49380# 8.08e-19
C8184 a_17408_49732# a_17408_49380# 0.0109f
C8185 XA2.XA4.MN0.D a_5960_49380# 0.154f
C8186 AVDD a_19928_43044# 0.00159f
C8187 D<1> a_18560_47620# 5.21e-19
C8188 D<5> a_8480_47268# 3.18e-19
C8189 a_12368_41636# a_13520_41636# 0.00133f
C8190 a_920_41636# XA0.XA1.XA1.MN0.S 0.0694f
C8191 SARP li_9184_30036# 0.00103f
C8192 XA0.XA4.MN0.G a_n232_47268# 0.157f
C8193 XA6.XA1.XA5.MN2.G a_14888_43748# 0.0732f
C8194 XA0.XA4.MN0.D a_n232_45860# 2.24e-19
C8195 AVDD a_18560_40580# 0.00125f
C8196 D<7> XA1.XA1.XA5.MN1.D 0.00185f
C8197 XA0.XA6.MP0.G a_920_44804# 5.5e-19
C8198 XA20.XA10.MN1.D XA20.XA9.MP0.D 2.14f
C8199 AVDD a_n232_52196# 0.00154f
C8200 a_n232_40228# a_920_40228# 0.00133f
C8201 XA4.XA4.MN0.G a_8480_44100# 2.84e-19
C8202 XA3.XA4.MN0.G a_9848_44100# 2.84e-19
C8203 VREF a_17408_43396# 3.39e-19
C8204 D<5> a_8480_41636# 6.49e-19
C8205 a_920_46212# a_920_45860# 0.0109f
C8206 XA4.XA3.MN0.G a_9848_45508# 0.104f
C8207 XA8.XA7.MP0.G XA8.XA1.XA1.MP2.D 0.0736f
C8208 XA3.XA1.XA5.MN2.G a_5960_41284# 0.0175f
C8209 D<1> a_18560_41988# 6.49e-19
C8210 AVDD a_11000_50084# 0.358f
C8211 XA3.XA9.MN1.G XA4.XA7.MP0.D 0.00108f
C8212 XA3.XA9.MN0.D XA3.XA7.MP0.D 0.00986f
C8213 CK_SAMPLE XA2.XA6.MN0.D 0.0659f
C8214 a_5960_52196# a_7328_52196# 8.89e-19
C8215 XA0.XA9.MN0.D a_n232_51844# 0.00176f
C8216 XA0.XA9.MN1.G a_920_51844# 6.57e-19
C8217 a_2288_52900# XA2.XA1.XA5.MN2.G 1.06e-19
C8218 XA7.XA9.MN0.D a_18560_52196# 0.0492f
C8219 XA7.XA9.MN1.G a_19928_52196# 2.84e-19
C8220 a_13808_1038# a_14960_1038# 0.00133f
C8221 XB2.XA3.MN0.S a_13808_334# 5.76e-19
C8222 XA0.XA4.MN0.G a_n232_41636# 6.69e-20
C8223 XA1.XA1.XA5.MN2.D a_3440_43748# 0.00224f
C8224 XA20.XA2a.MN0.D a_22448_43396# 0.00175f
C8225 XA7.XA1.XA5.MN2.D XA7.XA1.XA5.MN1.D 0.0488f
C8226 a_17408_45156# EN 1.83e-19
C8227 XA5.XA6.MP0.G a_12368_39876# 0.00273f
C8228 XA20.XA3a.MN0.D a_13520_42340# 0.00552f
C8229 AVDD D<8> 2.47f
C8230 XA5.XA1.XA5.MN2.G a_11000_50788# 0.00548f
C8231 a_2288_51140# a_2288_50788# 0.0109f
C8232 XA20.XA9.MP0.D a_23600_49028# 0.00334f
C8233 a_21080_52548# VREF 0.00386f
C8234 XA0.XA7.MP0.D a_n232_50084# 7.44e-20
C8235 a_14888_51140# XA6.XA6.MN2.D 0.00176f
C8236 a_16040_51140# D<2> 0.0672f
C8237 XB1.XA3.MN1.D m3_7544_1364# 0.0137f
C8238 XB2.XA4.MP0.D m3_16544_2420# 0.0634f
C8239 XA20.XA2a.MN0.D a_21080_40932# 0.0679f
C8240 XA2.XA3.MN0.G a_4808_40228# 0.00369f
C8241 EN XA0.XA1.XA4.MN0.D 0.00345f
C8242 a_17408_50084# a_18560_50084# 0.00133f
C8243 a_4808_50084# a_4808_49732# 0.0109f
C8244 XA6.XA1.XA5.MN2.G a_12368_47972# 0.00363f
C8245 XA7.XA6.MN0.D a_18560_49732# 0.00176f
C8246 D<1> a_17408_48676# 0.00918f
C8247 AVDD a_14888_43748# 0.00125f
C8248 D<5> a_7328_48324# 0.0164f
C8249 D<8> li_14804_20208# 3.5e-20
C8250 XA2.XA3.MN0.G XDAC2.XC128b<2>.XRES16.B 3.2e-20
C8251 a_5960_42340# a_5960_41988# 0.0109f
C8252 a_5960_42692# XA2.XA1.XA1.MN0.S 6.76e-20
C8253 XA7.XA6.MP0.G XA20.XA2a.MN0.D 0.0784f
C8254 XA4.XA6.MP0.G a_9848_46212# 4.4e-19
C8255 XA2.XA1.XA5.MN2.G a_4808_44452# 5.11e-19
C8256 XA0.XA6.MP0.G a_n232_45860# 7.76e-20
C8257 XA6.XA4.MN0.D a_14888_47268# 0.0963f
C8258 VREF a_22448_47268# 0.00162f
C8259 AVDD a_2288_41284# 0.361f
C8260 a_11000_48324# a_12368_48324# 8.89e-19
C8261 XA8.XA7.MP0.G a_22448_44804# 6.64e-19
C8262 AVDD XA8.XA10.MP0.D 0.728f
C8263 XA5.XA12.MP0.G XA6.XA12.MP0.G 0.00217f
C8264 XA20.XA11.MN0.D a_23600_53252# 0.071f
C8265 DONE a_22448_53252# 0.00598f
C8266 XA6.XA11.MN1.G XA8.XA11.MN1.G 1.54e-19
C8267 XA1.XA12.MP0.G a_2288_53604# 0.0877f
C8268 XA2.XA11.MN1.G a_3440_53604# 0.00787f
C8269 XA2.XA1.XA1.MN0.D a_4808_40580# 0.035f
C8270 XA7.XA1.XA1.MP1.D a_17408_40932# 0.0465f
C8271 a_13520_46916# a_13520_46564# 0.0109f
C8272 XA6.XA4.MN0.G XA5.XA1.XA5.MN2.D 0.0024f
C8273 XA5.XA4.MN0.G XA6.XA1.XA5.MN2.D 0.0024f
C8274 XA3.XA6.MP0.G a_7328_43396# 5.5e-19
C8275 XA5.XA3.MN0.G XA6.XA3.MN0.G 0.0258f
C8276 XA5.XA1.XA5.MN2.G a_12368_42340# 1.97e-19
C8277 XA7.XA6.MP0.G XA7.XA1.XA2.MP0.D 0.0125f
C8278 XA0.XA11.MN1.G XB1.XA2.MN0.G 0.0721f
C8279 XA20.XA4.MN0.D a_23600_52548# 0.0529f
C8280 CK_SAMPLE D<7> 0.0524f
C8281 AVDD a_9848_50788# 0.00154f
C8282 DONE XA8.XA6.MN2.D 2.25e-19
C8283 XB2.XA1.MP0.D XB2.XA4.MP0.D 0.0044f
C8284 SAR_IP a_11000_2094# 0.0503f
C8285 SARN XDAC2.XC0.XRES1A.B 3.59f
C8286 XA20.XA3a.MN0.D a_21080_43044# 0.00406f
C8287 XA4.XA1.XA5.MN2.D a_11000_44804# 0.156f
C8288 a_2288_45156# a_2288_44804# 0.0109f
C8289 a_14888_45156# a_16040_45156# 0.00133f
C8290 D<4> a_11000_39876# 7.76e-20
C8291 AVDD a_12368_47972# 0.356f
C8292 a_14888_51492# XA7.XA1.XA5.MN2.G 0.0674f
C8293 a_7328_53252# VREF 0.00267f
C8294 XA20.XA9.MP0.D a_23600_50084# 0.00614f
C8295 XDAC1.X16ab.XRES1B.B XDAC1.X16ab.XRES4.B 0.428f
C8296 XA20.XA2a.MN0.D XA1.XA1.XA1.MN0.S 0.137f
C8297 VREF CK_SAMPLE_BSSW 0.0297f
C8298 a_21080_43748# a_22448_43748# 8.89e-19
C8299 XA6.XA1.XA5.MP1.D XA6.XA1.XA5.MP0.D 0.0488f
C8300 XA1.XA1.XA5.MN1.D a_3440_43396# 0.00176f
C8301 EN a_8480_43396# 0.00238f
C8302 XA20.XA3a.MN0.D a_19928_40580# 0.0658f
C8303 a_18560_50436# XA7.XA6.MN0.D 0.00176f
C8304 XA5.XA1.XA5.MN2.G a_11000_49028# 0.00363f
C8305 AVDD a_n232_44452# 0.00125f
C8306 D<4> XA1.XA4.MN0.D 0.0609f
C8307 XA0.XA6.MP0.G XA6.XA6.MP0.G 0.0914f
C8308 XA1.XA6.MP0.G XA5.XA6.MP0.G 0.0592f
C8309 a_4808_50436# a_4808_50084# 0.0109f
C8310 XA2.XA6.MP0.G XA4.XA6.MP0.G 0.0287f
C8311 XDAC1.XC64a<0>.XRES8.B XDAC1.XC64a<0>.XRES16.B 0.0904f
C8312 li_9184_10992# li_9184_10380# 0.00271f
C8313 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC1.XRES1B.B 0.00444f
C8314 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES1A.B 0.0197f
C8315 XA1.XA1.XA2.MP0.D a_2288_41284# 1.07e-19
C8316 XA4.XA1.XA4.MN1.D a_9848_42340# 0.00176f
C8317 a_22448_42692# a_23600_42692# 0.00133f
C8318 D<8> XDAC1.XC0.XRES1A.B 9.7e-20
C8319 EN a_7328_40932# 0.00564f
C8320 a_4808_49028# a_4808_48676# 0.0109f
C8321 XA8.XA7.MP0.G a_21080_45860# 0.00363f
C8322 XA2.XA1.XA5.MN2.G a_4808_45508# 9.01e-20
C8323 AVDD a_11000_42340# 0.361f
C8324 VREF a_21080_48324# 0.0536f
C8325 D<5> a_8480_46212# 0.0141f
C8326 a_8480_54308# a_8480_53956# 0.0109f
C8327 a_21080_54308# a_22448_54308# 8.89e-19
C8328 AVDD XA4.XA11.MN1.G 1.04f
C8329 XA8.XA1.XA1.MN0.S a_21080_41284# 0.0964f
C8330 a_8480_41284# a_9848_41284# 8.89e-19
C8331 XA3.XA1.XA1.MN0.S XA3.XA1.XA1.MN0.D 0.0743f
C8332 XA3.XA1.XA1.MP2.D XA3.XA1.XA1.MP1.D 0.0488f
C8333 SARP XDAC1.XC128b<2>.XRES1A.B 3.59f
C8334 XA0.XA4.MN0.D a_n232_44804# 9.25e-20
C8335 XA6.XA6.MP0.G a_14888_44100# 7.76e-20
C8336 XA0.XA7.MP0.G XA0.XA1.XA4.MN1.D 7.2e-19
C8337 D<2> XA6.XA1.XA5.MP0.D 7.42e-19
C8338 AVDD XB2.XA1.MP0.D 0.433f
C8339 XA20.XA3a.MN0.D XA1.XA3.MN0.G 0.219f
C8340 XA1.XA4.MN0.G XA20.XA2a.MN0.D 0.00833f
C8341 XA0.XA4.MN0.G a_n232_46212# 0.0149f
C8342 XA7.XA4.MN0.G a_17408_46564# 3.46e-19
C8343 a_n232_47268# a_n232_46916# 0.0109f
C8344 D<6> a_5960_43396# 7.76e-20
C8345 AVDD a_16040_51492# 0.387f
C8346 XA5.XA11.MN1.G a_11000_52196# 4.29e-19
C8347 a_3440_52900# a_4808_52900# 8.89e-19
C8348 a_18560_39876# a_19928_39876# 8.89e-19
C8349 a_19928_45860# a_19928_45508# 0.0109f
C8350 XA3.XA3.MN0.G a_9848_44452# 6.55e-19
C8351 XA5.XA4.MN0.G XA5.XA1.XA5.MN0.D 0.0198f
C8352 D<6> a_4808_40932# 5.24e-19
C8353 XA7.XA1.XA5.MN2.G a_16040_40580# 0.0506f
C8354 SARN XB2.XA4.MP0.D 1.53f
C8355 XA2.XA4.MN0.D XA2.XA1.XA4.MN0.D 8.13e-19
C8356 XA20.XA3a.MN0.D a_16040_43748# 0.00106f
C8357 AVDD a_9848_49028# 0.00154f
C8358 XA6.XA7.MP0.D XA6.XA8.MP0.D 0.124f
C8359 a_2288_51844# XA1.XA8.MP0.D 0.0215f
C8360 a_13520_51844# a_14888_51844# 8.89e-19
C8361 XA1.XA7.MP0.D a_3440_51492# 0.126f
C8362 CK_SAMPLE XA5.XA4.MN0.D 0.0364f
C8363 XA3.XA9.MN1.G a_9848_51140# 2.84e-19
C8364 XA8.XA9.MN1.G XA8.XA1.XA5.MN2.G 4.35e-19
C8365 EN XA0.XA1.XA5.MP1.D 0.0545f
C8366 XA20.XA3a.MN0.D a_3440_41284# 0.00649f
C8367 XA20.XA2a.MN0.D XA5.XA1.XA4.MP0.D 0.0255f
C8368 XA2.XA1.XA5.MN2.D a_5960_43044# 1.88e-19
C8369 D<8> a_n232_41988# 0.00335f
C8370 XA20.XA9.MP0.D XA20.XA3a.MN0.D 0.058f
C8371 D<6> XA2.XA6.MP0.D 0.0323f
C8372 AVDD a_n232_45508# 0.00131f
C8373 a_16040_50788# a_17408_50788# 8.89e-19
C8374 XA5.XA1.XA5.MN2.G a_11000_50084# 0.00366f
C8375 a_2288_43044# a_2288_42692# 0.0109f
C8376 a_13520_43044# XA5.XA1.XA4.MN1.D 0.00176f
C8377 XA6.XA1.XA2.MP0.D XA6.XA1.XA4.MP0.D 4.34e-19
C8378 EN a_13520_41636# 1.25e-19
C8379 D<1> a_17408_47620# 0.0147f
C8380 XA3.XA1.XA5.MN2.G XA2.XA3.MN0.G 0.12f
C8381 XA2.XA4.MN0.D a_4808_49380# 0.155f
C8382 VREF a_7328_49380# 0.0171f
C8383 AVDD a_18560_43044# 0.00125f
C8384 D<5> a_7328_47268# 0.0148f
C8385 XA7.XA4.MN0.D XA8.XA4.MN0.D 0.00869f
C8386 a_12368_41988# XA5.XA1.XA1.MN0.S 3.8e-19
C8387 a_n232_41636# XA0.XA1.XA1.MN0.S 0.0674f
C8388 a_5960_47972# a_5960_47620# 0.0109f
C8389 XA6.XA4.MN0.G a_16040_47620# 0.155f
C8390 XA5.XA1.XA5.MN2.G a_14888_43748# 7.1e-20
C8391 XA6.XA1.XA5.MN2.G a_13520_43748# 2.66e-19
C8392 D<3> a_13520_44100# 6.49e-19
C8393 XA20.XA9.MP0.D a_23600_42340# 0.0674f
C8394 XA4.XA6.MP0.G a_11000_45156# 5.5e-19
C8395 XA6.XA4.MN0.D a_14888_46212# 1.1e-19
C8396 VREF a_22448_46212# 0.00165f
C8397 AVDD a_17408_40580# 0.381f
C8398 a_18560_47972# a_19928_47972# 8.89e-19
C8399 D<7> XA1.XA1.XA5.MP1.D 7.43e-19
C8400 D<6> EN 0.0613f
C8401 XA0.XA6.MP0.G a_n232_44804# 7.76e-20
C8402 XA20.XA10.MN1.D XA8.XA10.MP0.D 0.00217f
C8403 a_4808_53604# XA2.XA10.MP0.D 1.17e-19
C8404 a_16040_53604# a_16040_53252# 0.0109f
C8405 AVDD SARN 0.139f
C8406 a_12368_40580# a_12368_40228# 0.0109f
C8407 XA3.XA4.MN0.G a_8480_44100# 0.0164f
C8408 VREF a_16040_43396# 3.39e-19
C8409 XA0.XA11.MN1.G CK_SAMPLE_BSSW 4.96f
C8410 D<5> a_7328_41636# 7.77e-20
C8411 a_12368_46212# a_13520_46212# 0.00133f
C8412 XA3.XA3.MN0.G a_9848_45508# 7.98e-19
C8413 XA8.XA7.MP0.G XA8.XA1.XA1.MN0.S 0.305f
C8414 XA3.XA1.XA5.MN2.G a_4808_41284# 0.00527f
C8415 D<1> a_17408_41988# 7.77e-20
C8416 AVDD a_9848_50084# 0.00144f
C8417 XA3.XA9.MN1.G XA3.XA7.MP0.D 0.274f
C8418 CK_SAMPLE XA2.XA6.MP0.G 0.046f
C8419 XA5.XA10.MP0.G XA5.XA8.MP0.D 0.0434f
C8420 XA0.XA9.MN1.G a_n232_51844# 0.0164f
C8421 XA7.XA9.MN1.G a_18560_52196# 0.0878f
C8422 a_9560_1038# a_9560_686# 0.0109f
C8423 a_5960_44452# a_7328_44452# 8.89e-19
C8424 XA1.XA1.XA5.MN2.D a_2288_43748# 0.00388f
C8425 XA7.XA1.XA5.MN2.D XA7.XA1.XA5.MP1.D 0.0488f
C8426 XA6.XA4.MN0.G a_16040_41988# 5.1e-20
C8427 a_19928_44804# a_19928_44452# 0.0109f
C8428 a_16040_45156# EN 1.83e-19
C8429 SARN li_14804_20208# 0.00103f
C8430 XA5.XA6.MP0.G a_11000_39876# 1.28e-19
C8431 XA4.XA9.MN1.G a_11000_49732# 0.0215f
C8432 XA20.XA9.MP0.D a_22448_49028# 0.0714f
C8433 AVDD a_23600_46916# 0.00154f
C8434 XA5.XA1.XA5.MN2.G a_9848_50788# 1.87e-19
C8435 SARN XA20.XA3.MN0.D 0.422f
C8436 XB1.XA3.MN1.D m3_7472_1364# 0.0137f
C8437 XB2.XA4.MP0.D m3_16472_2420# 0.106f
C8438 li_14804_21432# li_14804_20820# 0.00271f
C8439 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128a<1>.XRES1B.B 0.00444f
C8440 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128b<2>.XRES16.B 0.0904f
C8441 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES1A.B 0.0197f
C8442 XA0.XA6.MP0.G XDAC2.XC32a<0>.XRES8.B 2.23e-21
C8443 XA20.XA2a.MN0.D a_19928_40932# 0.0718f
C8444 XA3.XA1.XA5.MN0.D a_8480_43044# 0.00176f
C8445 XA7.XA1.XA5.MN0.D a_18560_43396# 0.0474f
C8446 a_5960_43396# a_7328_43396# 8.89e-19
C8447 XA1.XA3.MN0.G a_4808_40228# 4.4e-20
C8448 XA2.XA3.MN0.G a_3440_40228# 4.21e-19
C8449 XA5.XA6.MP0.D VREF 0.0115f
C8450 XA6.XA1.XA5.MN2.G a_11000_47972# 7.1e-20
C8451 XA5.XA1.XA5.MN2.G a_12368_47972# 7.1e-20
C8452 AVDD a_13520_43748# 0.00125f
C8453 XA4.XA6.MP0.G XA4.XA4.MN0.D 0.76f
C8454 a_17408_42340# a_18560_42340# 0.00133f
C8455 XA7.XA1.XA4.MP0.D a_17408_41988# 0.00176f
C8456 XA2.XA1.XA5.MN2.G a_3440_44452# 1.86e-19
C8457 XA6.XA4.MN0.D a_13520_47268# 4.76e-20
C8458 XA5.XA4.MN0.D a_14888_47268# 4.76e-20
C8459 VREF a_21080_47268# 0.0188f
C8460 XA20.XA3.MN0.D a_23600_46916# 0.0275f
C8461 AVDD a_920_41284# 0.361f
C8462 a_23600_48676# a_23600_48324# 0.0109f
C8463 a_14888_48676# XA6.XA4.MN0.G 1.34e-19
C8464 XA8.XA7.MP0.G a_21080_44804# 0.00486f
C8465 AVDD XA7.XA10.MP0.D 0.727f
C8466 DONE a_21080_53252# 0.0015f
C8467 XA20.XA11.MN0.D a_22448_53252# 0.0658f
C8468 XA6.XA11.MN1.G XA6.XA12.MP0.G 0.214f
C8469 a_14888_53956# a_14888_53604# 0.0109f
C8470 XA2.XA11.MN1.G a_2288_53604# 0.00979f
C8471 XA1.XA1.XA1.MN0.S a_3440_39876# 2.54e-19
C8472 XA6.XA1.XA1.MN0.S a_16040_40228# 0.0313f
C8473 a_4808_40932# a_5960_40932# 0.00133f
C8474 SARP li_9184_9768# 0.00103f
C8475 D<8> a_920_46564# 0.155f
C8476 XA0.XA4.MN0.G a_920_45156# 5.54e-19
C8477 XA5.XA4.MN0.G XA5.XA1.XA5.MN2.D 0.135f
C8478 XA5.XA1.XA5.MN2.G a_11000_42340# 0.00442f
C8479 XA0.XA11.MN1.G a_9560_3502# 0.0379f
C8480 XA2.XA4.MN0.D XA2.XA1.XA5.MP1.D 9.69e-19
C8481 XA20.XA4.MN0.D a_22448_52548# 2.16e-19
C8482 a_9848_52548# a_11000_52548# 0.00133f
C8483 CK_SAMPLE XA0.XA6.MP2.D 3.06e-19
C8484 AVDD a_8480_50788# 0.00154f
C8485 DONE D<0> 0.00681f
C8486 XA2.XA10.MP0.G XA2.XA9.MN0.D 0.106f
C8487 SAR_IN XB2.XA4.MP0.D 0.00603f
C8488 SAR_IP a_9560_2094# 0.00157f
C8489 a_13808_2446# a_14960_2446# 0.00133f
C8490 a_9560_2446# XB1.XA4.MN0.D 0.00176f
C8491 XB2.XA1.MP0.D XB2.XA4.MN0.D 0.0109f
C8492 XA20.XA3a.MN0.D a_19928_43044# 0.0839f
C8493 XA4.XA1.XA5.MN2.D a_9848_44804# 0.153f
C8494 XA8.XA4.MN0.G XA8.XA1.XA4.MP1.D 0.0488f
C8495 XA2.XA4.MN0.G a_5960_42692# 0.00224f
C8496 XA7.XA3.MN0.G a_18560_43748# 2.78e-19
C8497 D<4> a_9848_39876# 0.00212f
C8498 SARN a_23600_50788# 0.088f
C8499 AVDD a_11000_47972# 0.356f
C8500 a_4808_51492# a_4808_51140# 0.0109f
C8501 XA4.XA9.MN1.G a_11000_50436# 7.76e-19
C8502 a_22448_51492# a_23600_51492# 0.00133f
C8503 a_5960_53252# VREF 0.00292f
C8504 XA20.XA2a.MN0.D XA0.XA1.XA1.MP2.D 0.0102f
C8505 EN a_7328_43396# 0.162f
C8506 XA20.XA3a.MN0.D a_18560_40580# 0.0674f
C8507 AVDD SARP 0.16f
C8508 D<4> VREF 1.3f
C8509 D<5> XA3.XA4.MN0.D 7.46f
C8510 XA8.XA1.XA4.MP1.D XA8.XA1.XA4.MP0.D 0.0488f
C8511 a_9848_42692# XA4.XA1.XA4.MN0.D 0.00176f
C8512 XA2.XA3.MN0.G XDAC2.XC0.XRES16.B 3.2e-20
C8513 D<8> li_14804_30648# 0.00508f
C8514 EN a_5960_40932# 0.00564f
C8515 a_16040_49028# a_17408_49028# 8.89e-19
C8516 D<1> a_18560_46564# 0.0551f
C8517 XA2.XA1.XA5.MN2.G a_3440_45508# 2.31e-19
C8518 AVDD a_9848_42340# 0.00125f
C8519 XA5.XA4.MN0.D a_13520_48324# 0.0997f
C8520 D<5> a_7328_46212# 0.0202f
C8521 AVDD XA2.XA12.MP0.G 0.709f
C8522 XA8.XA1.XA1.MN0.S a_19928_41284# 0.0658f
C8523 XA3.XA1.XA1.MN0.S XA3.XA1.XA1.MP1.D 0.0615f
C8524 XA20.XA3.MN0.D SARP 0.511f
C8525 XA3.XA6.MP0.G EN 0.065f
C8526 D<2> XA6.XA1.XA5.MN0.D 0.00188f
C8527 AVDD SAR_IN 0.0864f
C8528 XA20.XA3a.MN0.D D<8> 0.207f
C8529 XA0.XA4.MN0.G XA20.XA2a.MN0.D 0.00823f
C8530 a_11000_47268# a_12368_47268# 8.89e-19
C8531 D<6> a_4808_43396# 6.49e-19
C8532 XA7.XA1.XA5.MN2.G a_16040_43044# 0.00551f
C8533 CK_SAMPLE a_9848_51844# 1.64e-19
C8534 AVDD a_14888_51492# 0.00166f
C8535 XA20.XA10.MN1.D SARN 0.869f
C8536 a_22448_53252# a_22448_52900# 0.0109f
C8537 XA5.XA10.MP0.D a_13520_52900# 0.13f
C8538 a_9848_53604# XA4.XA9.MN1.G 7.36e-20
C8539 a_5960_45508# a_7328_45508# 8.89e-19
C8540 XA3.XA3.MN0.G a_8480_44452# 0.0963f
C8541 XA5.XA4.MN0.G XA5.XA1.XA5.MP0.D 0.00138f
C8542 SARN XB2.XA4.MN0.D 1.57e-19
C8543 XA7.XA1.XA5.MN2.G a_14888_40580# 9.75e-19
C8544 XA6.XA1.XA5.MN2.G a_16040_40580# 5.68e-19
C8545 XA20.XA3a.MN0.D a_14888_43748# 0.00218f
C8546 XA7.XA9.MN1.G XA8.XA7.MP0.G 4.35e-19
C8547 AVDD a_8480_49028# 0.00154f
C8548 XA1.XA7.MP0.D a_2288_51492# 0.0877f
C8549 CK_SAMPLE XA4.XA4.MN0.D 0.0364f
C8550 XA3.XA9.MN1.G a_8480_51140# 0.0469f
C8551 a_2288_52196# XA2.XA1.XA5.MN2.G 3.39e-19
C8552 XDAC1.XC0.XRES8.B XDAC1.XC0.XRES1A.B 0.0228f
C8553 XDAC1.XC0.XRES2.B XDAC1.XC0.XRES16.B 0.457f
C8554 EN XA0.XA1.XA5.MN1.D 0.0259f
C8555 SARN XDAC2.XC64a<0>.XRES16.B 55.3f
C8556 XA20.XA2a.MN0.D XA4.XA1.XA4.MP0.D 0.0251f
C8557 XA2.XA1.XA5.MN2.D a_4808_43044# 5.1e-20
C8558 XA0.XA6.MP2.G li_9184_25524# 3.5e-20
C8559 a_12368_44100# XA5.XA1.XA5.MP1.D 0.00176f
C8560 a_920_44100# a_920_43748# 0.0109f
C8561 a_3440_50788# a_3440_50436# 0.0109f
C8562 XA20.XA9.MP0.D a_23600_47972# 0.073f
C8563 D<6> XA2.XA6.MN0.D 0.00148f
C8564 XA6.XA6.MP2.D a_16040_50436# 0.00176f
C8565 AVDD a_23600_45860# 0.00154f
C8566 XA20.XA10.MN1.D a_23600_46916# 0.00423f
C8567 SARN a_23600_49028# 0.156f
C8568 a_22448_51844# VREF 0.00104f
C8569 XDAC1.XC128a<1>.XRES2.B XDAC1.XC32a<0>.XRES2.B 1.67e-19
C8570 li_9184_16116# li_9184_15696# 0.00411f
C8571 XA0.XA1.XA4.MN1.D XA0.XA1.XA4.MP1.D 0.00918f
C8572 XA2.XA1.XA2.MP0.D a_5960_42340# 2.54e-19
C8573 XA6.XA1.XA2.MP0.D XA6.XA1.XA4.MN0.D 0.056f
C8574 XA0.XA4.MN0.D XDAC1.XC32a<0>.XRES8.B 2.23e-21
C8575 EN a_12368_41636# 0.00649f
C8576 XA3.XA1.XA5.MN2.G XA1.XA3.MN0.G 1.07e-19
C8577 a_16040_49732# a_16040_49380# 0.0109f
C8578 VREF a_5960_49380# 0.0171f
C8579 XA2.XA1.XA5.MN2.G XA2.XA3.MN0.G 0.326f
C8580 AVDD a_17408_43044# 0.381f
C8581 a_11000_41636# a_12368_41636# 8.89e-19
C8582 SARP XDAC1.XC0.XRES1A.B 3.59f
C8583 XA6.XA4.MN0.G a_14888_47620# 0.154f
C8584 XA6.XA1.XA5.MN2.G a_12368_43748# 0.00442f
C8585 XA5.XA1.XA5.MN2.G a_13520_43748# 0.0749f
C8586 D<3> a_12368_44100# 7.77e-20
C8587 XA4.XA6.MP0.G a_9848_45156# 7.76e-20
C8588 XA20.XA3.MN0.D a_23600_45860# 0.0275f
C8589 VREF a_21080_46212# 0.067f
C8590 AVDD a_16040_40580# 0.381f
C8591 XA8.XA12.MP0.G XA8.XA10.MP0.D 0.0632f
C8592 XA3.XA12.MP0.G a_8480_52900# 0.00258f
C8593 XA4.XA11.MN1.G a_9848_52900# 7.39e-19
C8594 AVDD XA8.XA9.MN0.D 4.25e-19
C8595 XA3.XA4.MN0.G a_7328_44100# 6.11e-19
C8596 XA2.XA1.XA5.MN2.G a_4808_41284# 0.0044f
C8597 XA5.XA6.MP0.G a_13520_42692# 7.76e-20
C8598 a_n232_46212# a_n232_45860# 0.0109f
C8599 XA1.XA6.MP0.G XA1.XA1.XA4.MN0.D 6.07e-19
C8600 XA3.XA3.MN0.G a_8480_45508# 0.109f
C8601 XA8.XA1.XA5.MN2.G XA8.XA1.XA1.MN0.S 0.0308f
C8602 AVDD a_8480_50084# 0.00144f
C8603 a_4808_52196# a_5960_52196# 0.00133f
C8604 CK_SAMPLE XA1.XA6.MN0.D 0.0676f
C8605 a_920_52900# XA0.XA7.MP0.G 1.06e-19
C8606 XA7.XA9.MN1.G a_17408_52196# 0.0665f
C8607 a_9560_1390# CK_SAMPLE_BSSW 2.9e-19
C8608 a_12368_1038# a_13808_1038# 8e-19
C8609 XB2.XA0.MP0.D a_14960_n18# 0.00102f
C8610 XA20.XA2a.MN0.D a_19928_43396# 7.39e-20
C8611 XA6.XA4.MN0.G a_14888_41988# 1.74e-19
C8612 a_14888_45156# EN 4.58e-19
C8613 XA4.XA9.MN1.G a_9848_49732# 0.00119f
C8614 XA20.XA9.MP0.D a_21080_49028# 5.7e-20
C8615 AVDD a_22448_46916# 0.363f
C8616 a_920_51140# a_920_50788# 0.0109f
C8617 D<7> D<6> 1.33f
C8618 XA0.XA6.MP2.G D<5> 0.185f
C8619 SARN a_23600_50084# 0.0882f
C8620 XB1.XA3.MN1.D m3_n1960_2244# 0.0634f
C8621 XB2.XA4.MP0.D m3_26048_3300# 0.0273f
C8622 XA20.XA2a.MN0.D a_18560_40932# 0.0733f
C8623 XA7.XA1.XA5.MN0.D a_17408_43396# 2.16e-19
C8624 XA7.XA1.XA5.MP0.D a_18560_43396# 2.16e-19
C8625 XA1.XA3.MN0.G a_3440_40228# 0.00307f
C8626 EN a_22448_42692# 5.7e-20
C8627 XA5.XA6.MP0.G VREF 0.568f
C8628 XA5.XA1.XA5.MN2.G a_11000_47972# 0.00363f
C8629 XA20.XA10.MN1.D SARP 0.423f
C8630 XA1.XA6.MP0.G a_3440_49380# 0.0547f
C8631 AVDD a_12368_43748# 0.357f
C8632 XA4.XA6.MP0.G XA3.XA4.MN0.D 0.00194f
C8633 XA7.XA6.MP0.G a_18560_49732# 0.00239f
C8634 XA7.XA6.MP0.D a_17408_49732# 0.00176f
C8635 a_3440_50084# a_3440_49732# 0.0109f
C8636 a_16040_50084# a_17408_50084# 8.89e-19
C8637 a_4808_42340# a_4808_41988# 0.0109f
C8638 D<8> XDAC2.XC128b<2>.XRES16.B 3.84e-19
C8639 AVDD a_n232_41284# 0.00125f
C8640 D<5> a_8480_45156# 7.77e-19
C8641 VREF a_19928_47268# 1.19e-19
C8642 XA5.XA4.MN0.D a_13520_47268# 0.0963f
C8643 a_9848_48324# a_11000_48324# 0.00133f
C8644 XA8.XA7.MP0.G a_19928_44804# 1.86e-19
C8645 XA2.XA1.XA5.MN2.G a_2288_44452# 0.00486f
C8646 XA0.XA7.MP0.G a_3440_44452# 5.11e-19
C8647 XA0.XA12.MP0.D a_3440_53604# 0.0726f
C8648 DONE a_19928_53252# 5.02e-20
C8649 XA6.XA11.MN1.G XA7.XA11.MN1.G 0.0251f
C8650 XA2.XA11.MN1.G a_920_53604# 9.49e-20
C8651 AVDD XA6.XA10.MP0.D 0.728f
C8652 XA1.XA1.XA1.MN0.S a_2288_39876# 2.54e-19
C8653 XA6.XA1.XA1.MN0.S a_14888_40228# 0.0215f
C8654 XA1.XA1.XA1.MN0.D a_3440_40580# 0.035f
C8655 XA6.XA1.XA1.MP1.D a_16040_40932# 0.0465f
C8656 a_12368_46916# a_12368_46564# 0.0109f
C8657 D<8> a_n232_46564# 0.156f
C8658 XA0.XA4.MN0.G a_n232_45156# 0.00865f
C8659 XA4.XA3.MN0.G XA5.XA3.MN0.G 0.00869f
C8660 XA5.XA1.XA5.MN2.G a_9848_42340# 3.12e-19
C8661 XA4.XA1.XA5.MN2.G a_11000_42340# 1.97e-19
C8662 VREF XA3.XA1.XA5.MP1.D 0.00623f
C8663 XA2.XA4.MN0.D XA2.XA1.XA5.MN1.D 9.9e-19
C8664 CK_SAMPLE XA0.XA6.MN2.D 0.0389f
C8665 AVDD a_7328_50788# 0.363f
C8666 XA2.XA10.MP0.G XA2.XA9.MN1.G 0.202f
C8667 XB1.XA1.MN0.D a_9560_2094# 4.63e-19
C8668 a_11000_2446# XB1.M1.G 1.61e-19
C8669 XB2.XA1.MP0.D XB2.M1.G 0.129f
C8670 XB2.XA1.MN0.D XB2.XA4.MP0.D 0.0122f
C8671 SARN li_14804_30648# 0.00103f
C8672 XA20.XA3a.MN0.D a_18560_43044# 0.0905f
C8673 a_13520_45156# a_14888_45156# 8.89e-19
C8674 a_920_45156# a_920_44804# 0.0109f
C8675 XA6.XA6.MP0.G XA6.XA1.XA1.MN0.D 0.00159f
C8676 XA8.XA4.MN0.G XA8.XA1.XA4.MN1.D 0.0642f
C8677 XA2.XA4.MN0.G a_4808_42692# 0.0049f
C8678 D<4> a_8480_39876# 8.39e-20
C8679 a_7328_51844# D<5> 1.25e-19
C8680 XA6.XA7.MP0.D D<2> 2.65e-19
C8681 SARN a_22448_50788# 5.88e-19
C8682 AVDD a_9848_47972# 0.00125f
C8683 a_13520_51492# XA6.XA1.XA5.MN2.G 0.0658f
C8684 XA4.XA9.MN1.G a_9848_50436# 0.01f
C8685 li_14804_26556# li_14804_26136# 0.00411f
C8686 XDAC2.XC64b<1>.XRES2.B XDAC2.X16ab.XRES2.B 1.67e-19
C8687 a_5960_43748# XA2.XA1.XA5.MP0.D 0.00176f
C8688 a_19928_43748# a_21080_43748# 0.00133f
C8689 XA6.XA1.XA5.MN1.D XA6.XA1.XA5.MN0.D 0.0488f
C8690 XA6.XA1.XA5.MP1.D XA6.XA1.XA2.MP0.D 6.52e-20
C8691 XA20.XA2a.MN0.D XA0.XA1.XA1.MN0.S 0.137f
C8692 XA3.XA3.MN0.G a_9848_41284# 7.98e-19
C8693 XA1.XA1.XA5.MP1.D a_2288_43396# 0.00176f
C8694 EN a_5960_43396# 0.162f
C8695 XA20.XA3a.MN0.D a_17408_40580# 0.0658f
C8696 SARN XA20.XA3a.MN0.D 2.71e-19
C8697 AVDD a_23600_44804# 0.00159f
C8698 D<4> XA0.XA4.MN0.D 0.0525f
C8699 D<5> XA2.XA4.MN0.D 3.83f
C8700 a_18560_50436# XA7.XA6.MP0.G 3.02e-20
C8701 a_17408_50436# XA7.XA6.MP0.D 0.00176f
C8702 a_3440_50436# a_3440_50084# 0.0109f
C8703 XA20.XA10.MN1.D a_23600_45860# 0.00423f
C8704 XDAC2.XC64a<0>.XRES8.B XDAC2.XC64a<0>.XRES2.B 0.44f
C8705 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES1A.B 0.00438f
C8706 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES16.B 0.0483f
C8707 XA8.XA1.XA2.MP0.D a_21080_41636# 0.00224f
C8708 XA3.XA1.XA4.MN1.D a_8480_42340# 0.00176f
C8709 a_21080_42692# a_22448_42692# 8.89e-19
C8710 XA1.XA3.MN0.G XDAC2.XC0.XRES16.B 5.78e-20
C8711 D<3> XA20.XA2a.MN0.D 0.0858f
C8712 a_3440_49028# a_3440_48676# 0.0109f
C8713 D<1> a_17408_46564# 0.0695f
C8714 XA2.XA1.XA5.MN2.G a_2288_45508# 0.00595f
C8715 XA0.XA7.MP0.G a_3440_45508# 9.01e-20
C8716 AVDD a_8480_42340# 0.00125f
C8717 XA5.XA4.MN0.D a_12368_48324# 0.0682f
C8718 a_19928_54308# a_21080_54308# 0.00133f
C8719 AVDD XA3.XA11.MN1.G 1.89f
C8720 a_7328_54308# a_7328_53956# 0.0109f
C8721 XA20.XA12.MP0.G a_22448_53956# 0.00201f
C8722 XA20.XA12.MP0.D a_23600_53956# 0.0661f
C8723 a_7328_41284# a_8480_41284# 0.00133f
C8724 SARP li_9184_20208# 0.00103f
C8725 AVDD XB2.XA1.MN0.D 0.514f
C8726 VREF a_22448_45156# 0.0016f
C8727 XA20.XA3.MN0.D a_23600_44804# 0.0287f
C8728 SARN a_23600_42340# 0.00204f
C8729 D<2> XA6.XA1.XA2.MP0.D 0.0153f
C8730 XA20.XA3a.MN0.D a_23600_46916# 0.0533f
C8731 XA6.XA4.MN0.G a_16040_46564# 3.46e-19
C8732 a_23600_47620# a_23600_47268# 0.0109f
C8733 XA7.XA1.XA5.MN2.G a_14888_43044# 2.31e-19
C8734 CK_SAMPLE a_8480_51844# 2.08e-19
C8735 AVDD a_13520_51492# 0.00166f
C8736 XA5.XA10.MP0.D a_12368_52900# 0.0877f
C8737 a_2288_52900# a_3440_52900# 0.00133f
C8738 a_17408_39876# a_18560_39876# 0.00133f
C8739 D<3> XA5.XA1.XA1.MN0.D 0.0166f
C8740 a_18560_45860# a_18560_45508# 0.0109f
C8741 XA3.XA3.MN0.G a_7328_44452# 0.055f
C8742 XA5.XA4.MN0.G XA5.XA1.XA2.MP0.D 0.206f
C8743 SARN XB2.M1.G 0.285f
C8744 XA6.XA1.XA5.MN2.G a_14888_40580# 0.083f
C8745 XA1.XA4.MN0.D XA1.XA1.XA4.MN0.D 8.11e-19
C8746 XA20.XA3a.MN0.D a_13520_43748# 0.00228f
C8747 XA7.XA9.MN1.G XA8.XA1.XA5.MN2.G 0.0494f
C8748 AVDD a_7328_49028# 0.356f
C8749 XA5.XA7.MP0.D XA5.XA8.MP0.D 0.124f
C8750 a_920_51844# XA0.XA8.MP0.D 0.0215f
C8751 a_12368_51844# a_13520_51844# 0.00133f
C8752 CK_SAMPLE XA3.XA4.MN0.D 0.0364f
C8753 a_2288_53956# VREF 0.00396f
C8754 XA3.XA9.MN1.G a_7328_51140# 0.0222f
C8755 XA8.XA1.XA5.MN2.D a_21080_43396# 4.58e-19
C8756 XA20.XA2a.MN0.D XA4.XA1.XA4.MN0.D 0.0375f
C8757 D<6> XA2.XA6.MP0.G 0.468f
C8758 D<4> XA0.XA6.MP0.G 0.0861f
C8759 XA20.XA9.MP0.D a_22448_47972# 0.0658f
C8760 AVDD a_22448_45860# 0.403f
C8761 XA20.XA10.MN1.D a_22448_46916# 1.89e-19
C8762 a_14888_50788# a_16040_50788# 0.00133f
C8763 D<5> XA1.XA6.MP0.G 0.0629f
C8764 a_21080_51844# VREF 0.0037f
C8765 a_920_43044# a_920_42692# 0.0109f
C8766 a_12368_43044# XA5.XA1.XA4.MP1.D 0.00176f
C8767 XA2.XA1.XA2.MP0.D a_4808_42340# 0.095f
C8768 EN a_11000_41636# 0.00649f
C8769 AVDD a_16040_43044# 0.381f
C8770 VREF a_4808_49380# 8.08e-19
C8771 XA7.XA6.MP0.G a_18560_48676# 0.0651f
C8772 XA0.XA7.MP0.G XA2.XA3.MN0.G 0.0241f
C8773 XA2.XA1.XA5.MN2.G XA1.XA3.MN0.G 0.222f
C8774 XA6.XA4.MN0.D XA7.XA4.MN0.D 0.00869f
C8775 XA1.XA4.MN0.D a_3440_49380# 0.155f
C8776 XA3.XA6.MP0.G a_8480_48324# 0.00295f
C8777 a_23600_41988# a_23600_41636# 0.0109f
C8778 a_4808_47972# a_4808_47620# 0.0109f
C8779 XA7.XA6.MP0.G XA7.XA1.XA5.MN2.D 0.0325f
C8780 XA5.XA4.MN0.D a_13520_46212# 1.1e-19
C8781 VREF a_19928_46212# 7.12e-19
C8782 AVDD a_14888_40580# 0.00125f
C8783 a_17408_47972# a_18560_47972# 0.00133f
C8784 XA3.XA12.MP0.G a_7328_52900# 1.28e-19
C8785 XA4.XA11.MN1.G a_8480_52900# 0.00295f
C8786 a_3440_53604# XA1.XA10.MP0.D 1.17e-19
C8787 a_14888_53604# a_14888_53252# 0.0109f
C8788 XA1.XA11.MP0.D a_2288_53252# 0.0494f
C8789 AVDD XA8.XA9.MN1.G 0.926f
C8790 a_11000_40580# a_11000_40228# 0.0109f
C8791 XA5.XA6.MP0.G a_12368_42692# 5.5e-19
C8792 XA20.XA3a.MN0.D SARP 9.59e-20
C8793 a_11000_46212# a_12368_46212# 8.89e-19
C8794 XA1.XA6.MP0.G XA1.XA1.XA4.MP0.D 9.97e-19
C8795 XA3.XA3.MN0.G a_7328_45508# 0.0682f
C8796 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MP2.D 0.0739f
C8797 XA7.XA1.XA5.MN2.G XA8.XA1.XA1.MN0.S 5.21e-19
C8798 XA2.XA1.XA5.MN2.G a_3440_41284# 0.00733f
C8799 XA0.XA11.MN1.G a_13808_686# 0.00206f
C8800 AVDD a_7328_50084# 0.358f
C8801 XA2.XA9.MN0.D XA2.XA7.MP0.D 0.00986f
C8802 CK_SAMPLE XA1.XA6.MP0.D 0.0278f
C8803 DONE XA8.XA6.MP0.D 4.24e-20
C8804 XA4.XA10.MP0.G XA4.XA8.MP0.D 0.0434f
C8805 XA0.XA10.MP0.G a_n232_51492# 6.8e-20
C8806 XA20.XA4.MN0.D a_23600_51844# 0.056f
C8807 a_8408_1038# a_8408_686# 0.0109f
C8808 XB2.XA0.MP0.D a_13808_n18# 6.02e-19
C8809 a_4808_44452# a_5960_44452# 0.00133f
C8810 XA20.XA2a.MN0.D a_18560_43396# 4.8e-20
C8811 XA0.XA1.XA5.MN2.D a_920_43748# 0.00388f
C8812 XA6.XA1.XA5.MN2.D XA6.XA1.XA5.MP1.D 0.0488f
C8813 XA8.XA3.MN0.G a_19928_43044# 3.62e-20
C8814 a_13520_45156# EN 4.58e-19
C8815 a_18560_44804# a_18560_44452# 0.0109f
C8816 XA4.XA6.MP0.G a_12368_39876# 5.53e-19
C8817 XA3.XA4.MN0.D a_8480_40932# 9.24e-20
C8818 SARN XDAC2.XC128b<2>.XRES16.B 55.3f
C8819 XA20.XA3a.MN0.D a_9848_42340# 0.00547f
C8820 AVDD a_21080_46916# 0.359f
C8821 XA4.XA1.XA5.MN2.G a_8480_50788# 1.87e-19
C8822 D<7> XA1.XA6.MN2.D 1.59e-19
C8823 a_17408_52548# VREF 0.00396f
C8824 SARN a_22448_50084# 5.34e-19
C8825 a_13520_51140# XA5.XA6.MN2.D 0.00176f
C8826 XB1.XA3.MN1.D m3_n2104_2244# 0.17f
C8827 XB2.XA4.MP0.D m3_25976_3300# 0.0137f
C8828 li_9184_21432# li_9184_20820# 0.00271f
C8829 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128a<1>.XRES1B.B 0.00444f
C8830 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128b<2>.XRES16.B 0.0904f
C8831 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES1A.B 0.0197f
C8832 XA0.XA6.MP0.G li_14804_15084# 1.85e-20
C8833 XA20.XA2a.MN0.D a_17408_40932# 0.0662f
C8834 SARP a_23600_42340# 0.0892f
C8835 XA3.XA1.XA2.MP0.D a_8480_43044# 0.0292f
C8836 XA3.XA1.XA5.MP0.D a_7328_43044# 0.00176f
C8837 XA7.XA1.XA5.MP0.D a_17408_43396# 0.049f
C8838 a_4808_43396# a_5960_43396# 0.00133f
C8839 XA7.XA1.XA2.MP0.D a_18560_43396# 0.0961f
C8840 EN a_21080_42692# 0.159f
C8841 XA4.XA6.MP0.D VREF 0.0115f
C8842 XA20.XA10.MN1.D a_23600_44804# 0.005f
C8843 XA1.XA6.MP0.G a_2288_49380# 0.0781f
C8844 AVDD a_11000_43748# 0.357f
C8845 XA7.XA6.MP0.G a_17408_49732# 0.099f
C8846 a_16040_42340# a_17408_42340# 8.89e-19
C8847 XA6.XA1.XA4.MP0.D a_16040_41988# 0.00176f
C8848 XA7.XA1.XA2.MP0.D a_17408_40932# 4.25e-20
C8849 SARP XB2.M1.G 0.0183f
C8850 AVDD XA8.XA1.XA1.MP2.D 0.127f
C8851 D<2> XA6.XA1.XA5.MN2.D 0.0347f
C8852 D<5> a_7328_45156# 6.68e-19
C8853 VREF a_18560_47268# 1.19e-19
C8854 XA5.XA4.MN0.D a_12368_47268# 0.0576f
C8855 XA6.XA6.MP0.G XA20.XA2a.MN0.D 0.0783f
C8856 a_22448_48676# a_22448_48324# 0.0109f
C8857 a_13520_48676# XA5.XA4.MN0.G 1.34e-19
C8858 XA8.XA1.XA5.MN2.G a_19928_44804# 1.95e-19
C8859 XA0.XA7.MP0.G a_2288_44452# 7.1e-20
C8860 XA2.XA1.XA5.MN2.G a_920_44452# 7.1e-20
C8861 XA6.XA11.MN1.G XA5.XA12.MP0.G 0.391f
C8862 XA0.XA12.MP0.D a_2288_53604# 0.073f
C8863 XA0.XA12.MP0.G a_920_53604# 0.0893f
C8864 a_13520_53956# a_13520_53604# 0.0109f
C8865 XA5.XA11.MN1.G XA6.XA12.MP0.G 0.00122f
C8866 AVDD XA5.XA10.MP0.D 0.727f
C8867 XA1.XA1.XA1.MN0.D a_2288_40580# 8.3e-19
C8868 XA6.XA1.XA1.MN0.D a_16040_40932# 8.29e-20
C8869 a_3440_40932# a_4808_40932# 8.89e-19
C8870 SARP XDAC1.XC64a<0>.XRES16.B 55.3f
C8871 XA4.XA4.MN0.G XA4.XA1.XA5.MN2.D 0.135f
C8872 XA0.XA6.MP2.G XA0.XA1.XA4.MP0.D 6.08e-19
C8873 XA4.XA1.XA5.MN2.G a_9848_42340# 0.00568f
C8874 D<4> a_11000_42692# 7.76e-20
C8875 XA0.XA11.MN1.G a_9560_3854# 0.00283f
C8876 VREF XA2.XA1.XA5.MP1.D 0.00623f
C8877 XA20.XA3a.MN0.D a_23600_45860# 8.07e-19
C8878 a_8480_52548# a_9848_52548# 8.89e-19
C8879 XA8.XA10.MP0.G a_21080_52548# 0.07f
C8880 CK_SAMPLE XA0.XA6.MP2.G 0.0523f
C8881 AVDD a_5960_50788# 0.363f
C8882 XB1.XA1.MP0.D a_9560_2094# 0.0738f
C8883 a_12368_2446# a_13808_2446# 8e-19
C8884 a_9560_2446# XB1.M1.G 0.0339f
C8885 a_8408_2446# XB1.XA4.MP0.D 0.00977f
C8886 SAR_IN XB2.M1.G 0.682f
C8887 XA2.XA6.MP0.G a_5960_40932# 4.24e-19
C8888 XA20.XA3a.MN0.D a_17408_43044# 0.00877f
C8889 XA3.XA1.XA5.MN2.D a_8480_44804# 0.153f
C8890 D<8> XA0.XA1.XA2.MP0.D 0.0351f
C8891 AVDD a_8480_47972# 0.00125f
C8892 a_3440_51492# a_3440_51140# 0.0109f
C8893 a_12368_51492# XA6.XA1.XA5.MN2.G 0.0714f
C8894 a_21080_51492# a_22448_51492# 8.89e-19
C8895 XA6.XA1.XA5.MN1.D XA6.XA1.XA2.MP0.D 0.0102f
C8896 XA3.XA3.MN0.G a_8480_41284# 0.00342f
C8897 EN a_4808_43396# 0.00238f
C8898 XA20.XA3a.MN0.D a_16040_40580# 0.0674f
C8899 SARN a_23600_47972# 0.00206f
C8900 AVDD a_22448_44804# 0.366f
C8901 XA1.XA6.MP0.G XA4.XA6.MP0.G 0.0596f
C8902 XA0.XA6.MP2.G a_920_49380# 0.00891f
C8903 XA2.XA6.MP0.G XA3.XA6.MP0.G 1.9f
C8904 D<5> XA1.XA4.MN0.D 0.267f
C8905 XA3.XA6.MP2.D VREF 5.13e-19
C8906 a_17408_50436# XA7.XA6.MP0.G 0.0678f
C8907 D<2> a_16040_49732# 0.0109f
C8908 XA20.XA10.MN1.D a_22448_45860# 2.14e-19
C8909 XA0.XA6.MP0.G XA5.XA6.MP0.G 0.0759f
C8910 XA8.XA1.XA4.MN1.D XA8.XA1.XA4.MN0.D 0.0488f
C8911 XA4.XA1.XA2.MP0.D XA4.XA1.XA1.MN0.S 2.11e-19
C8912 XA8.XA1.XA2.MP0.D a_19928_41636# 0.00316f
C8913 a_8480_42692# XA3.XA1.XA4.MN0.D 0.00176f
C8914 D<8> XDAC2.XC0.XRES16.B 0.0333f
C8915 a_14888_49028# a_16040_49028# 0.00133f
C8916 XA3.XA6.MP0.G a_8480_47268# 1.38e-19
C8917 XA20.XA9.MP0.D a_23600_43748# 0.00334f
C8918 XA0.XA7.MP0.G a_2288_45508# 7.1e-20
C8919 XA2.XA1.XA5.MN2.G a_920_45508# 7.1e-20
C8920 AVDD a_7328_42340# 0.361f
C8921 VREF a_17408_48324# 0.0536f
C8922 XA7.XA6.MP0.G a_18560_47620# 4.4e-19
C8923 XA20.XA12.MP0.G a_21080_53956# 0.047f
C8924 XA20.XA12.MP0.D a_22448_53956# 0.0986f
C8925 AVDD XA1.XA12.MP0.G 0.706f
C8926 XA2.XA1.XA1.MP2.D XA2.XA1.XA1.MP1.D 0.0488f
C8927 AVDD SAR_IP 0.0864f
C8928 VREF a_21080_45156# 0.0192f
C8929 XA20.XA3a.MN0.D a_22448_46916# 0.0608f
C8930 XA6.XA4.MN0.G a_14888_46564# 0.0155f
C8931 a_9848_47268# a_11000_47268# 0.00133f
C8932 XA6.XA1.XA5.MN2.G a_14888_43044# 0.0748f
C8933 XA1.XA6.MP0.G XA1.XA1.XA5.MN1.D 7.41e-19
C8934 a_21080_53252# a_21080_52900# 0.0109f
C8935 AVDD a_12368_51492# 0.387f
C8936 a_4808_45508# a_5960_45508# 0.00133f
C8937 a_7328_45860# XA3.XA1.XA5.MN2.D 3.12e-20
C8938 XA3.XA6.MP0.G a_8480_41636# 7.76e-20
C8939 XA5.XA1.XA5.MN2.G a_14888_40580# 7.1e-20
C8940 XA6.XA1.XA5.MN2.G a_13520_40580# 0.00564f
C8941 XA7.XA6.MP0.G a_18560_41988# 7.76e-20
C8942 XA1.XA4.MN0.D XA1.XA1.XA4.MP0.D 7.97e-19
C8943 XA20.XA3a.MN0.D a_12368_43748# 0.00106f
C8944 AVDD a_5960_49028# 0.356f
C8945 a_n232_51844# XA0.XA8.MP0.D 0.0215f
C8946 XA0.XA7.MP0.D a_920_51492# 0.0893f
C8947 CK_SAMPLE XA2.XA4.MN0.D 0.0364f
C8948 a_920_53956# VREF 0.00366f
C8949 a_920_52196# XA0.XA7.MP0.G 3.39e-19
C8950 XDAC2.XC0.XRES8.B XDAC2.XC0.XRES16.B 0.0904f
C8951 li_14804_31872# li_14804_31260# 0.00271f
C8952 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES1A.B 0.0197f
C8953 XDAC2.XC0.XRES1B.B XDAC2.XC64b<1>.XRES1B.B 0.00444f
C8954 XA20.XA3a.MN0.D a_n232_41284# 0.00643f
C8955 SARN li_14804_10380# 0.00103f
C8956 XA8.XA1.XA5.MN2.D a_19928_43396# 1.28e-19
C8957 XA20.XA2a.MN0.D XA3.XA1.XA4.MN0.D 0.0409f
C8958 XA1.XA1.XA5.MN2.D a_3440_43044# 5.1e-20
C8959 a_n232_44452# XA0.XA1.XA2.MP0.D 5.16e-20
C8960 XA0.XA6.MP2.G XDAC1.X16ab.XRES4.B 4.06e-21
C8961 a_11000_44100# XA4.XA1.XA5.MP1.D 0.00176f
C8962 a_n232_44100# a_n232_43748# 0.0109f
C8963 a_2288_50788# a_2288_50436# 0.0109f
C8964 D<2> a_16040_50436# 0.0879f
C8965 XA6.XA6.MN2.D a_14888_50436# 0.00176f
C8966 a_16040_51140# XA6.XA6.MP0.G 6.76e-20
C8967 AVDD a_21080_45860# 0.356f
C8968 XDAC2.XC128a<1>.XRES1A.B XDAC2.XC32a<0>.XRES1B.B 0.617f
C8969 EN a_9848_41636# 1.25e-19
C8970 XA0.XA4.MN0.D li_9184_15084# 1.85e-20
C8971 XA7.XA6.MP0.G a_17408_48676# 0.0881f
C8972 XA2.XA1.XA5.MN2.G D<8> 6.95e-19
C8973 XA0.XA7.MP0.G XA1.XA3.MN0.G 0.229f
C8974 AVDD a_14888_43044# 0.00125f
C8975 XA8.XA1.XA5.MN2.G a_17408_46916# 0.00455f
C8976 a_14888_49732# a_14888_49380# 0.0109f
C8977 XA1.XA4.MN0.D a_2288_49380# 0.154f
C8978 VREF a_3440_49380# 8.08e-19
C8979 XA3.XA6.MP0.G a_7328_48324# 0.00417f
C8980 a_11000_41988# XA4.XA1.XA1.MN0.S 3.8e-19
C8981 a_9848_41636# a_11000_41636# 0.00133f
C8982 SARP li_9184_30648# 0.00103f
C8983 XA5.XA4.MN0.G a_13520_47620# 0.154f
C8984 XA5.XA1.XA5.MN2.G a_11000_43748# 0.00442f
C8985 VREF a_18560_46212# 7.12e-19
C8986 AVDD a_13520_40580# 0.00125f
C8987 D<7> EN 0.0614f
C8988 XA20.XA3.MN6.D a_23600_45508# 0.154f
C8989 XA7.XA12.MP0.G XA7.XA10.MP0.D 0.0632f
C8990 XA8.XA11.MN1.G XA8.XA10.MP0.D 0.0625f
C8991 AVDD XA7.XA9.MN0.D 4.25e-19
C8992 XA4.XA11.MN1.G a_7328_52900# 1.34e-19
C8993 a_22448_40580# a_23600_40580# 0.00133f
C8994 XA2.XA4.MN0.G a_5960_44100# 6.11e-19
C8995 VREF a_12368_43396# 3.39e-19
C8996 XA3.XA4.MN0.D a_8480_43396# 9.24e-20
C8997 XA20.XA2a.MN0.D a_23600_46212# 0.0528f
C8998 XA8.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.S 0.301f
C8999 XA0.XA7.MP0.G a_3440_41284# 0.00392f
C9000 XA2.XA1.XA5.MN2.G a_2288_41284# 0.0169f
C9001 XA0.XA11.MN1.G a_12368_686# 0.00139f
C9002 AVDD a_5960_50084# 0.358f
C9003 XA2.XA9.MN1.G XA2.XA7.MP0.D 0.274f
C9004 a_3440_52196# a_4808_52196# 8.89e-19
C9005 CK_SAMPLE XA1.XA6.MP0.G 0.0463f
C9006 DONE XA8.XA6.MN0.D 4.24e-20
C9007 XA20.XA4.MN0.D a_22448_51844# 2.43e-19
C9008 a_11000_1038# a_12368_1038# 8.89e-19
C9009 XB1.XA3.MN1.D a_9560_334# 9.07e-19
C9010 XB2.XA3.MN1.D CK_SAMPLE_BSSW 0.0531f
C9011 XA0.XA1.XA5.MN2.D a_n232_43748# 0.00224f
C9012 XA6.XA1.XA5.MN2.D XA6.XA1.XA5.MN1.D 0.0488f
C9013 XA5.XA4.MN0.G a_13520_41988# 1.74e-19
C9014 a_12368_45156# EN 1.83e-19
C9015 XA4.XA6.MP0.G a_11000_39876# 0.00322f
C9016 XA3.XA4.MN0.D a_7328_40932# 9.15e-20
C9017 XA20.XA3a.MN0.D a_8480_42340# 0.00552f
C9018 AVDD a_19928_46916# 0.00166f
C9019 XA4.XA1.XA5.MN2.G a_7328_50788# 0.00548f
C9020 a_n232_51140# a_n232_50788# 0.0109f
C9021 D<7> XA1.XA6.MP2.D 0.0399f
C9022 a_16040_52548# VREF 0.00396f
C9023 XB1.XA3.MN1.D m3_7544_2420# 0.0137f
C9024 XB2.XA4.MP0.D m3_16544_3476# 0.0634f
C9025 XA20.XA2a.MN0.D a_16040_40932# 0.0678f
C9026 SARP a_22448_42340# 5.54e-19
C9027 XA3.XA1.XA2.MP0.D a_7328_43044# 3.59e-19
C9028 XA20.XA10.MN1.D a_22448_44804# 1.69e-19
C9029 D<6> a_5960_48324# 0.0164f
C9030 AVDD a_9848_43748# 0.00125f
C9031 D<2> a_16040_48676# 0.00918f
C9032 a_2288_50084# a_2288_49732# 0.0109f
C9033 a_14888_50084# a_16040_50084# 0.00133f
C9034 a_3440_42340# a_3440_41988# 0.0109f
C9035 SARP XB1.XA4.MN0.D 1.57e-19
C9036 D<8> li_14804_20820# 3.5e-20
C9037 AVDD XA8.XA1.XA1.MN0.S 1.05f
C9038 VREF a_17408_47268# 0.0191f
C9039 XA3.XA6.MP0.G a_8480_46212# 7.76e-20
C9040 a_8480_48324# a_9848_48324# 8.89e-19
C9041 XA8.XA1.XA5.MN2.G a_18560_44804# 1.86e-19
C9042 XA0.XA7.MP0.G a_920_44452# 0.00486f
C9043 XA0.XA12.MP0.D a_920_53604# 0.0124f
C9044 XA0.XA12.MP0.G a_n232_53604# 0.1f
C9045 XA4.XA12.MP0.G XA5.XA12.MP0.G 0.00217f
C9046 AVDD XA4.XA10.MP0.D 0.728f
C9047 XA1.XA1.XA1.MP1.D a_2288_40580# 0.00176f
C9048 XA6.XA1.XA1.MN0.D a_14888_40932# 0.0535f
C9049 a_11000_46916# a_11000_46564# 0.0109f
C9050 XA4.XA4.MN0.G XA3.XA1.XA5.MN2.D 0.0024f
C9051 XA3.XA4.MN0.G XA4.XA1.XA5.MN2.D 0.0024f
C9052 XA6.XA6.MP0.G XA6.XA1.XA5.MP0.D 0.00121f
C9053 XA3.XA3.MN0.G XA4.XA3.MN0.G 0.0261f
C9054 XA0.XA6.MP2.G XA0.XA1.XA4.MN0.D 0.00144f
C9055 XA4.XA1.XA5.MN2.G a_8480_42340# 4.69e-19
C9056 D<4> a_9848_42692# 6.49e-19
C9057 XA2.XA6.MP0.G a_5960_43396# 5.5e-19
C9058 XA1.XA4.MN0.D XA1.XA1.XA5.MN1.D 9.89e-19
C9059 XA20.XA3a.MN0.D a_22448_45860# 0.00498f
C9060 a_14888_52900# XA6.XA9.MN1.G 0.00113f
C9061 XA8.XA10.MP0.G a_19928_52548# 0.128f
C9062 XA1.XA10.MP0.G XA1.XA9.MN0.D 0.106f
C9063 CK_SAMPLE a_23600_51140# 7.93e-19
C9064 AVDD a_4808_50788# 0.00154f
C9065 a_8408_2446# XB1.M1.G 0.0712f
C9066 XB2.XA1.MN0.D XB2.M1.G 0.0319f
C9067 XB1.XA1.MP0.D a_8408_2094# 2.01e-19
C9068 a_8408_3150# XB1.XA3.MN1.D 0.00238f
C9069 XA2.XA6.MP0.G a_4808_40932# 3.97e-20
C9070 SARN XDAC2.XC0.XRES16.B 55.3f
C9071 XA20.XA3a.MN0.D a_16040_43044# 0.00835f
C9072 a_12368_45156# a_13520_45156# 0.00133f
C9073 XA3.XA1.XA5.MN2.D a_7328_44804# 0.156f
C9074 a_n232_45156# a_n232_44804# 0.0109f
C9075 XA7.XA4.MN0.G XA7.XA1.XA4.MN1.D 0.0642f
C9076 XA1.XA4.MN0.G a_3440_42692# 0.0049f
C9077 AVDD a_7328_47972# 0.356f
C9078 a_2288_53252# VREF 0.00267f
C9079 li_9184_26556# li_9184_26136# 0.00411f
C9080 XDAC1.XC64b<1>.XRES2.B XDAC1.X16ab.XRES2.B 1.67e-19
C9081 a_4808_43748# XA2.XA1.XA5.MN0.D 0.00176f
C9082 a_18560_43748# a_19928_43748# 8.89e-19
C9083 XA20.XA2a.MN0.D a_22448_41636# 0.00207f
C9084 XA0.XA1.XA5.MP1.D a_920_43396# 0.00176f
C9085 EN a_3440_43396# 0.00238f
C9086 XA20.XA3a.MN0.D a_14888_40580# 0.0658f
C9087 AVDD a_21080_44804# 0.356f
C9088 XA0.XA6.MP2.G a_n232_49380# 5.91e-19
C9089 D<6> XA3.XA4.MN0.D 0.0317f
C9090 XA2.XA6.MP0.G XA2.XA6.MP0.D 0.0392f
C9091 D<5> VREF 1.3f
C9092 D<2> a_14888_49732# 7.01e-19
C9093 a_2288_50436# a_2288_50084# 0.0109f
C9094 XA4.XA1.XA5.MN2.G a_7328_49028# 0.00363f
C9095 XDAC2.XC64a<0>.XRES8.B li_14804_10992# 9.91e-20
C9096 XDAC1.XC64a<0>.XRES8.B XDAC1.XC64a<0>.XRES2.B 0.44f
C9097 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES1A.B 0.00438f
C9098 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES16.B 0.0483f
C9099 XA0.XA1.XA2.MP0.D a_920_41284# 1.07e-19
C9100 XA3.XA1.XA4.MP1.D a_7328_42340# 0.00176f
C9101 a_19928_42692# a_21080_42692# 0.00133f
C9102 D<8> XDAC1.XC0.XRES16.B 0.00155f
C9103 EN a_2288_40932# 0.00564f
C9104 XA8.XA1.XA5.MN2.G a_17408_45860# 0.00363f
C9105 a_2288_49028# a_2288_48676# 0.0109f
C9106 XA3.XA6.MP0.G a_7328_47268# 5.95e-19
C9107 XA20.XA9.MP0.D a_22448_43748# 0.072f
C9108 XA0.XA7.MP0.G a_920_45508# 0.00595f
C9109 AVDD a_5960_42340# 0.361f
C9110 VREF a_16040_48324# 0.0536f
C9111 XA4.XA4.MN0.D a_11000_48324# 0.0698f
C9112 XA7.XA6.MP0.G a_17408_47620# 6.35e-19
C9113 a_18560_54308# a_19928_54308# 8.89e-19
C9114 a_5960_54308# a_5960_53956# 0.0109f
C9115 XA20.XA12.MP0.G a_19928_53956# 0.0224f
C9116 AVDD XA2.XA11.MN1.G 1.04f
C9117 XA7.XA1.XA1.MN0.S a_18560_41284# 0.0674f
C9118 a_5960_41284# a_7328_41284# 8.89e-19
C9119 XA7.XA1.XA1.MP2.D a_17408_41284# 0.0465f
C9120 XA2.XA1.XA1.MN0.S XA2.XA1.XA1.MP1.D 0.0615f
C9121 SARP XDAC1.XC128b<2>.XRES16.B 55.3f
C9122 AVDD XB1.XA1.MN0.D 0.514f
C9123 XA20.XA3a.MN0.D a_21080_46916# 2.07e-19
C9124 XA2.XA6.MP0.G EN 0.0651f
C9125 XA5.XA6.MP0.G a_13520_44100# 7.76e-20
C9126 XA20.XA3a.MN0.G a_23600_44452# 8.29e-20
C9127 XA20.XA3.MN6.D a_22448_44452# 0.16f
C9128 XA5.XA4.MN0.G a_14888_46564# 2.2e-19
C9129 XA6.XA4.MN0.G a_13520_46564# 2.2e-19
C9130 a_22448_47620# a_22448_47268# 0.0109f
C9131 XA6.XA1.XA5.MN2.G a_13520_43044# 2.31e-19
C9132 XA1.XA6.MP0.G XA1.XA1.XA5.MP1.D 0.00121f
C9133 VREF a_19928_45156# 7.39e-19
C9134 XA8.XA12.MP0.G XA8.XA9.MN1.G 4.5e-19
C9135 XA4.XA11.MN1.G a_8480_52196# 1.84e-19
C9136 XA4.XA10.MP0.D a_11000_52900# 0.0893f
C9137 a_920_52900# a_2288_52900# 8.89e-19
C9138 AVDD a_11000_51492# 0.387f
C9139 a_16040_39876# a_17408_39876# 8.89e-19
C9140 XA20.XA2a.MN0.D XA20.XA2.MN1.D 0.103f
C9141 a_17408_45860# a_17408_45508# 0.0109f
C9142 D<7> a_3440_40932# 5.26e-19
C9143 XA2.XA3.MN0.G a_5960_44452# 0.055f
C9144 XA4.XA4.MN0.G XA4.XA1.XA5.MP0.D 0.00138f
C9145 XA3.XA6.MP0.G a_7328_41636# 5.5e-19
C9146 XA5.XA1.XA5.MN2.G a_13520_40580# 0.0806f
C9147 XA6.XA1.XA5.MN2.G a_12368_40580# 0.0431f
C9148 XA7.XA6.MP0.G a_17408_41988# 5.5e-19
C9149 XA20.XA3a.MN0.D a_11000_43748# 0.00106f
C9150 AVDD a_4808_49028# 0.00154f
C9151 XA4.XA7.MP0.D XA4.XA8.MP0.D 0.124f
C9152 a_11000_51844# a_12368_51844# 8.89e-19
C9153 XA0.XA7.MP0.D a_n232_51492# 0.124f
C9154 CK_SAMPLE XA1.XA4.MN0.D 0.0364f
C9155 XA20.XA2a.MN0.D XA3.XA1.XA4.MP0.D 0.0255f
C9156 XA1.XA1.XA5.MN2.D a_2288_43044# 1.88e-19
C9157 a_9848_44804# XA4.XA1.XA2.MP0.D 2.6e-20
C9158 D<2> a_14888_50436# 5.7e-19
C9159 AVDD a_19928_45860# 0.00129f
C9160 a_13520_50788# a_14888_50788# 8.89e-19
C9161 XA4.XA1.XA5.MN2.G a_7328_50084# 0.00366f
C9162 a_n232_43044# a_n232_42692# 0.0109f
C9163 a_11000_43044# XA4.XA1.XA4.MP1.D 0.00176f
C9164 EN a_8480_41636# 1.25e-19
C9165 XA0.XA7.MP0.G D<8> 0.12f
C9166 AVDD a_13520_43044# 0.00125f
C9167 D<2> a_16040_47620# 0.0147f
C9168 VREF a_2288_49380# 0.0171f
C9169 XA5.XA4.MN0.D XA6.XA4.MN0.D 0.00869f
C9170 D<6> a_5960_47268# 0.0148f
C9171 XA7.XA1.XA5.MN2.G a_17408_46916# 7.1e-20
C9172 XA8.XA1.XA5.MN2.G a_16040_46916# 7.1e-20
C9173 XA20.XA1.MN0.D a_23600_41284# 0.056f
C9174 a_22448_41988# a_22448_41636# 0.0109f
C9175 XA5.XA1.XA5.MN2.G a_9848_43748# 1.95e-19
C9176 XA5.XA4.MN0.G a_12368_47620# 0.155f
C9177 VREF a_17408_46212# 0.0671f
C9178 AVDD a_12368_40580# 0.381f
C9179 a_16040_47972# a_17408_47972# 8.89e-19
C9180 XA0.XA6.MP2.G XA0.XA1.XA5.MP1.D 7.42e-19
C9181 XA20.XA3.MN6.D a_22448_45508# 0.168f
C9182 a_3440_47972# a_3440_47620# 0.0109f
C9183 XA8.XA11.MN1.G XA7.XA10.MP0.D 0.0327f
C9184 AVDD XA7.XA9.MN1.G 0.93f
C9185 XA3.XA11.MN1.G a_8480_52900# 0.00208f
C9186 a_13520_53604# a_13520_53252# 0.0109f
C9187 XA0.XA11.MP0.D a_920_53252# 0.0494f
C9188 a_9848_40580# a_9848_40228# 0.0109f
C9189 D<2> a_16040_41988# 7.76e-20
C9190 XA20.XA3a.MN0.D a_22448_44804# 0.0044f
C9191 XA20.XA2a.MN0.D a_22448_46212# 0.0438f
C9192 a_9848_46212# a_11000_46212# 0.00133f
C9193 a_23600_46564# a_23600_46212# 0.0109f
C9194 XA2.XA3.MN0.G a_5960_45508# 0.0698f
C9195 D<6> a_5960_41636# 7.76e-20
C9196 XA7.XA1.XA5.MN2.G XA7.XA1.XA1.MN0.S 0.0916f
C9197 XA0.XA7.MP0.G a_2288_41284# 5.96e-19
C9198 XA0.XA11.MN1.G a_11000_686# 0.00139f
C9199 XA3.XA4.MN0.D a_7328_43396# 9.15e-20
C9200 VREF a_11000_43396# 3.39e-19
C9201 XA2.XA4.MN0.G a_4808_44100# 0.0164f
C9202 AVDD a_4808_50084# 0.00144f
C9203 XA2.XA9.MN1.G XA1.XA7.MP0.D 0.00108f
C9204 XA6.XA9.MN0.D a_14888_52196# 0.0492f
C9205 CK_SAMPLE XA0.XA6.MP0.D 0.0276f
C9206 DONE XA8.XA6.MP0.G 8.91e-20
C9207 XA3.XA10.MP0.G XA3.XA8.MP0.D 0.0434f
C9208 XA20.XA9.MP0.D a_23600_51492# 0.00339f
C9209 XA6.XA9.MN1.G a_16040_52196# 0.0681f
C9210 XB1.XA3.MN0.S a_9560_334# 5.76e-19
C9211 XB2.XA4.MP0.D m3_26048_132# 0.0273f
C9212 XB1.XA3.MN1.D a_8408_334# 0.00886f
C9213 XB2.XA3.MN0.S CK_SAMPLE_BSSW 0.00496f
C9214 XB2.XA3.MN1.D a_14960_686# 0.00656f
C9215 a_14960_1390# a_14960_1038# 0.0109f
C9216 a_3440_44452# a_4808_44452# 8.89e-19
C9217 XA7.XA3.MN0.G a_18560_43044# 3.62e-20
C9218 XA5.XA4.MN0.G a_12368_41988# 5.1e-20
C9219 a_11000_45156# EN 1.83e-19
C9220 a_17408_44804# a_17408_44452# 0.0109f
C9221 XA4.XA6.MP0.G a_9848_39876# 7.76e-20
C9222 SARN li_14804_20820# 0.00103f
C9223 XA0.XA6.MP2.G D<6> 0.00792f
C9224 AVDD a_18560_46916# 0.00131f
C9225 XA3.XA1.XA5.MN2.G a_7328_50788# 7.1e-20
C9226 XA4.XA1.XA5.MN2.G a_5960_50788# 7.1e-20
C9227 XA3.XA9.MN1.G a_8480_49732# 0.00119f
C9228 a_12368_51140# XA5.XA6.MP2.D 0.00176f
C9229 XB1.XA3.MN1.D m3_7472_2420# 0.0137f
C9230 XB2.XA4.MP0.D m3_16472_3476# 0.106f
C9231 XDAC2.XC128b<2>.XRES8.B XDAC2.XC128b<2>.XRES2.B 0.44f
C9232 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES16.B 0.0483f
C9233 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES1A.B 0.00438f
C9234 XA0.XA6.MP0.G XDAC2.XC32a<0>.XRES4.B 2.23e-21
C9235 XA20.XA2a.MN0.D a_14888_40932# 0.0717f
C9236 a_3440_43396# a_4808_43396# 8.89e-19
C9237 D<6> a_4808_48324# 6.53e-19
C9238 AVDD a_8480_43748# 0.00125f
C9239 XA3.XA6.MP0.G XA3.XA4.MN0.D 4.49f
C9240 D<2> a_14888_48676# 3.48e-19
C9241 XA4.XA6.MP0.G VREF 0.568f
C9242 XA6.XA6.MP0.D a_16040_49732# 0.00176f
C9243 li_14804_6288# li_14804_5676# 0.00271f
C9244 a_14888_42340# a_16040_42340# 0.00133f
C9245 XA6.XA1.XA4.MN0.D a_14888_41988# 0.00176f
C9246 a_2288_42692# XA1.XA1.XA1.MN0.S 6.76e-20
C9247 SARP XB1.XA4.MP0.D 1.54f
C9248 XA4.XA4.MN0.D a_11000_47268# 0.0576f
C9249 VREF a_16040_47268# 0.0191f
C9250 AVDD XA7.XA1.XA1.MP2.D 0.127f
C9251 SARN a_23600_43748# 0.0017f
C9252 XA3.XA6.MP0.G a_7328_46212# 5.5e-19
C9253 a_21080_48676# a_21080_48324# 0.0109f
C9254 XA8.XA1.XA5.MN2.G a_17408_44804# 0.00486f
C9255 XA7.XA1.XA5.MN2.G a_18560_44804# 1.95e-19
C9256 XA0.XA7.MP0.G a_n232_44452# 1.86e-19
C9257 XA7.XA6.MP0.G a_18560_46564# 5e-19
C9258 a_n232_53956# XA0.XA11.MN1.G 7.59e-19
C9259 XA0.XA12.MP0.D a_n232_53604# 0.00305f
C9260 a_12368_53956# a_12368_53604# 0.0109f
C9261 XA20.XA12.MP0.G a_21080_53252# 0.00144f
C9262 XA20.XA12.MP0.D a_22448_53252# 3.8e-19
C9263 XA5.XA11.MN1.G XA5.XA12.MP0.G 0.278f
C9264 XA4.XA12.MP0.G XA6.XA11.MN1.G 1.54e-19
C9265 AVDD XA3.XA10.MP0.D 0.727f
C9266 XA0.XA1.XA1.MN0.S a_920_39876# 2.54e-19
C9267 XA5.XA1.XA1.MN0.S a_13520_40228# 0.0215f
C9268 a_2288_40932# a_3440_40932# 0.00133f
C9269 SARP li_9184_10380# 0.00103f
C9270 XA4.XA1.XA5.MN2.G a_7328_42340# 0.00442f
C9271 XA3.XA1.XA5.MN2.G a_8480_42340# 0.00568f
C9272 XA3.XA4.MN0.G XA3.XA1.XA5.MN2.D 0.135f
C9273 XA6.XA6.MP0.G XA6.XA1.XA5.MN0.D 7.41e-19
C9274 XA2.XA6.MP0.G a_4808_43396# 7.76e-20
C9275 XA1.XA4.MN0.D XA1.XA1.XA5.MP1.D 9.71e-19
C9276 XA20.XA3a.MN0.D a_21080_45860# 3.15e-19
C9277 a_7328_52548# a_8480_52548# 0.00133f
C9278 XA1.XA10.MP0.G XA1.XA9.MN1.G 0.202f
C9279 CK_SAMPLE a_22448_51140# 0.00817f
C9280 AVDD a_3440_50788# 0.00154f
C9281 a_11000_2446# a_12368_2446# 8.89e-19
C9282 SAR_IP XB2.M1.G 4.38e-19
C9283 XA20.XA3a.MN0.D a_14888_43044# 0.0864f
C9284 D<5> a_8480_39876# 0.00173f
C9285 XA7.XA4.MN0.G XA7.XA1.XA4.MP1.D 0.0488f
C9286 XA1.XA4.MN0.G a_2288_42692# 0.00224f
C9287 XA6.XA3.MN0.G a_14888_43748# 2.78e-19
C9288 D<1> a_18560_40228# 2.88e-19
C9289 XA8.XA9.MN1.G a_21080_50788# 0.00281f
C9290 AVDD a_5960_47972# 0.356f
C9291 XA3.XA9.MN1.G a_8480_50436# 0.01f
C9292 a_2288_51492# a_2288_51140# 0.0109f
C9293 a_11000_51492# XA5.XA1.XA5.MN2.G 0.0699f
C9294 a_19928_51492# a_21080_51492# 0.00133f
C9295 a_920_53252# VREF 0.00292f
C9296 a_4808_43748# XA2.XA1.XA2.MP0.D 0.0702f
C9297 XA5.XA1.XA5.MN1.D XA5.XA1.XA5.MN0.D 0.0488f
C9298 XA20.XA2a.MN0.D a_21080_41636# 0.00245f
C9299 EN a_2288_43396# 0.162f
C9300 XA20.XA3a.MN0.D a_13520_40580# 0.0674f
C9301 AVDD a_19928_44804# 0.00154f
C9302 XA2.XA6.MP2.D VREF 5.13e-19
C9303 D<6> XA2.XA4.MN0.D 7.43f
C9304 D<5> XA0.XA4.MN0.D 0.455f
C9305 a_16040_50436# XA6.XA6.MP0.D 0.00176f
C9306 XA3.XA1.XA5.MN2.G a_7328_49028# 7.1e-20
C9307 XA4.XA1.XA5.MN2.G a_5960_49028# 7.1e-20
C9308 XA7.XA1.XA4.MN1.D XA7.XA1.XA4.MN0.D 0.0488f
C9309 a_7328_42692# XA3.XA1.XA4.MP0.D 0.00176f
C9310 D<8> li_14804_31260# 0.00508f
C9311 EN a_920_40932# 0.00581f
C9312 D<4> XA20.XA2a.MN0.D 0.0851f
C9313 XA8.XA1.XA5.MN2.G a_16040_45860# 7.1e-20
C9314 XA7.XA1.XA5.MN2.G a_17408_45860# 7.1e-20
C9315 D<6> a_5960_46212# 0.0202f
C9316 a_13520_49028# a_14888_49028# 8.89e-19
C9317 XA20.XA9.MP0.D a_21080_43748# 5.7e-20
C9318 XA0.XA7.MP0.G a_n232_45508# 2.31e-19
C9319 AVDD a_4808_42340# 0.00125f
C9320 XA4.XA4.MN0.D a_9848_48324# 0.0981f
C9321 AVDD XA0.XA12.MP0.G 0.709f
C9322 XA7.XA1.XA1.MN0.S a_17408_41284# 0.0948f
C9323 XA2.XA1.XA1.MN0.S XA2.XA1.XA1.MN0.D 0.0743f
C9324 AVDD XB1.XA1.MP0.D 0.433f
C9325 XA5.XA6.MP0.G a_12368_44100# 5.5e-19
C9326 XA20.XA3a.MN0.G a_22448_44452# 0.0142f
C9327 XA5.XA4.MN0.G a_13520_46564# 0.0155f
C9328 a_8480_47268# a_9848_47268# 8.89e-19
C9329 D<7> a_3440_43396# 6.49e-19
C9330 XA5.XA1.XA5.MN2.G a_13520_43044# 0.0732f
C9331 XA6.XA1.XA5.MN2.G a_12368_43044# 0.00551f
C9332 VREF a_18560_45156# 7.39e-19
C9333 a_19928_53252# a_19928_52900# 0.0109f
C9334 XA4.XA10.MP0.D a_9848_52900# 0.128f
C9335 AVDD a_9848_51492# 0.00166f
C9336 CK_SAMPLE a_4808_51844# 1.64e-19
C9337 XA20.XA2a.MN0.D a_23600_45156# 0.00668f
C9338 XA5.XA1.XA5.MN2.G a_12368_40580# 0.00417f
C9339 D<7> a_2288_40932# 4.18e-20
C9340 XA2.XA3.MN0.G a_4808_44452# 0.096f
C9341 XA4.XA4.MN0.G XA4.XA1.XA5.MN0.D 0.0198f
C9342 SARN XB1.M1.G 0.141f
C9343 XA20.XA3a.MN0.D a_9848_43748# 0.00218f
C9344 a_5960_45860# XA2.XA1.XA5.MN2.D 3.12e-20
C9345 a_3440_45508# a_4808_45508# 8.89e-19
C9346 XA6.XA9.MN1.G XA7.XA1.XA5.MN2.G 0.0494f
C9347 AVDD a_3440_49028# 0.00154f
C9348 CK_SAMPLE VREF 1.93f
C9349 XA2.XA9.MN1.G a_5960_51140# 0.0222f
C9350 XDAC1.XC0.XRES8.B XDAC1.XC0.XRES16.B 0.0904f
C9351 li_9184_31872# li_9184_31260# 0.00271f
C9352 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES1A.B 0.0197f
C9353 XDAC1.XC0.XRES1B.B XDAC1.XC64b<1>.XRES1B.B 0.00444f
C9354 SARN XDAC2.XC64a<0>.XRES2.B 6.99f
C9355 XA20.XA3a.MN0.D XA8.XA1.XA1.MN0.S 0.0673f
C9356 a_21080_44100# EN 0.0752f
C9357 a_22448_44100# a_23600_44100# 0.00133f
C9358 XA7.XA1.XA5.MN2.D a_18560_43396# 1.28e-19
C9359 XA20.XA2a.MN0.D XA2.XA1.XA4.MP0.D 0.0251f
C9360 a_19928_45156# XA8.XA1.XA2.MP0.D 1.56e-20
C9361 SARP a_23600_43748# 0.155f
C9362 XA0.XA6.MP2.G li_9184_26136# 3.5e-20
C9363 a_9848_44100# XA4.XA1.XA5.MN1.D 0.00176f
C9364 a_920_50788# a_920_50436# 0.0109f
C9365 D<5> XA0.XA6.MP0.G 0.0629f
C9366 D<6> XA1.XA6.MP0.G 0.0712f
C9367 AVDD a_18560_45860# 0.00125f
C9368 XA4.XA1.XA5.MN2.G a_5960_50084# 7.1e-20
C9369 XA3.XA1.XA5.MN2.G a_7328_50084# 7.1e-20
C9370 a_17408_51844# VREF 0.00396f
C9371 XDAC1.XC128a<1>.XRES1A.B XDAC1.XC32a<0>.XRES1B.B 0.617f
C9372 a_22448_43044# a_23600_43044# 0.00133f
C9373 XA5.XA1.XA2.MP0.D XA5.XA1.XA4.MN0.D 0.056f
C9374 EN a_7328_41636# 0.00649f
C9375 XA0.XA4.MN0.D XDAC1.XC32a<0>.XRES4.B 2.23e-21
C9376 a_13520_49732# a_13520_49380# 0.0109f
C9377 AVDD a_12368_43044# 0.381f
C9378 D<2> a_14888_47620# 5.21e-19
C9379 VREF a_920_49380# 0.0171f
C9380 D<6> a_4808_47268# 3.18e-19
C9381 XA7.XA1.XA5.MN2.G a_16040_46916# 0.00455f
C9382 XA20.XA1.MN0.D a_22448_41284# 2.67e-19
C9383 a_8480_41636# a_9848_41636# 8.89e-19
C9384 SARP XDAC1.XC0.XRES16.B 55.3f
C9385 XA3.XA6.MP0.G a_8480_45156# 7.76e-20
C9386 XA4.XA1.XA5.MN2.G a_9848_43748# 0.0732f
C9387 D<0> a_21080_44452# 1.06e-19
C9388 VREF a_16040_46212# 0.0671f
C9389 AVDD a_11000_40580# 0.381f
C9390 XA0.XA6.MP2.G XA0.XA1.XA5.MN1.D 0.00185f
C9391 D<4> a_11000_44100# 7.76e-20
C9392 XA20.XA3a.MN0.G a_22448_45508# 0.0277f
C9393 AVDD XA6.XA9.MN0.D 4.25e-19
C9394 XA2.XA12.MP0.G a_5960_52900# 1.28e-19
C9395 XA3.XA11.MN1.G a_7328_52900# 0.00273f
C9396 XA0.XA11.MN1.G a_920_53252# 0.0674f
C9397 a_21080_40580# a_22448_40580# 8.89e-19
C9398 D<2> a_14888_41988# 6.49e-19
C9399 XA2.XA3.MN0.G a_4808_45508# 0.107f
C9400 D<6> a_4808_41636# 6.49e-19
C9401 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MP2.D 0.0736f
C9402 XA8.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S 3.84e-21
C9403 XA0.XA7.MP0.G a_920_41284# 0.0175f
C9404 XA0.XA11.MN1.G a_9560_686# 0.00206f
C9405 XA1.XA4.MN0.G a_4808_44100# 2.84e-19
C9406 XA2.XA4.MN0.G a_3440_44100# 2.84e-19
C9407 XA8.XA4.MN0.G a_21080_44452# 5.54e-19
C9408 CK_SAMPLE XA0.XA6.MN0.D 0.0659f
C9409 XA6.XA9.MN1.G a_14888_52196# 0.0862f
C9410 a_2288_52196# a_3440_52196# 0.00133f
C9411 a_19928_52548# XA8.XA7.MP0.D 5.16e-20
C9412 XA1.XA9.MN0.D XA1.XA7.MP0.D 0.00986f
C9413 XA8.XA10.MP0.G a_21080_51844# 0.00224f
C9414 XA1.XA9.MN1.G XA2.XA7.MP0.D 0.00108f
C9415 AVDD a_3440_50084# 0.00144f
C9416 XB2.XA4.MP0.D m3_25976_132# 0.0137f
C9417 XB1.XA3.MN1.D CK_SAMPLE_BSSW 0.046f
C9418 XB2.XA3.MN0.S a_14960_686# 0.0215f
C9419 XB2.XA3.MN1.D a_13808_686# 4.45e-19
C9420 a_9560_1038# a_11000_1038# 8e-19
C9421 XA3.XA6.MP0.G a_12368_39876# 2.67e-19
C9422 XA20.XA2a.MN0.D a_14888_43396# 7.39e-20
C9423 a_9848_45156# EN 4.58e-19
C9424 XA2.XA4.MN0.D a_5960_40932# 9.14e-20
C9425 XA5.XA1.XA5.MN2.D XA5.XA1.XA5.MN1.D 0.0488f
C9426 XA8.XA7.MP0.G XA8.XA6.MP2.D 0.00313f
C9427 AVDD a_17408_46916# 0.359f
C9428 XA3.XA1.XA5.MN2.G a_5960_50788# 0.00548f
C9429 XA3.XA9.MN1.G a_7328_49732# 0.0215f
C9430 XA8.XA9.MN1.G a_21080_50084# 0.00281f
C9431 a_12368_51140# D<3> 0.0688f
C9432 XB1.XA3.MN1.D m3_n1960_3300# 0.0634f
C9433 XB2.XA4.MP0.D m3_26048_4356# 0.0273f
C9434 XA20.XA2a.MN0.D a_13520_40932# 0.0733f
C9435 XA2.XA1.XA5.MP0.D a_5960_43044# 0.00176f
C9436 XA6.XA1.XA5.MP0.D a_16040_43396# 0.049f
C9437 D<8> a_n232_40228# 0.00369f
C9438 EN a_17408_42692# 0.159f
C9439 XA4.XA1.XA5.MN2.G a_7328_47972# 0.00363f
C9440 AVDD a_7328_43748# 0.357f
C9441 XA3.XA6.MP0.G XA2.XA4.MN0.D 2.8e-19
C9442 a_920_50084# a_920_49732# 0.0109f
C9443 a_13520_50084# a_14888_50084# 8.89e-19
C9444 a_2288_42340# a_2288_41988# 0.0109f
C9445 SARP XB1.M1.G 0.228f
C9446 D<8> XDAC2.XC128b<2>.XRES2.B 4.06e-21
C9447 VREF a_14888_47268# 1.19e-19
C9448 XA4.XA4.MN0.D a_9848_47268# 0.0963f
C9449 AVDD XA7.XA1.XA1.MN0.S 1.03f
C9450 XA5.XA6.MP0.G XA20.XA2a.MN0.D 0.0784f
C9451 D<0> a_21080_45508# 0.00428f
C9452 a_7328_48324# a_8480_48324# 0.00133f
C9453 XA7.XA1.XA5.MN2.G a_17408_44804# 7.1e-20
C9454 XA8.XA1.XA5.MN2.G a_16040_44804# 7.1e-20
C9455 XA7.XA6.MP0.G a_17408_46564# 5.5e-19
C9456 XA5.XA11.MN1.G XA6.XA11.MN1.G 0.271f
C9457 AVDD XA2.XA10.MP0.D 0.728f
C9458 XA0.XA1.XA1.MN0.S a_n232_39876# 2.54e-19
C9459 XA5.XA1.XA1.MN0.S a_12368_40228# 0.0313f
C9460 XA0.XA1.XA1.MP1.D a_920_40580# 0.00176f
C9461 XA5.XA1.XA1.MN0.D a_13520_40932# 0.0535f
C9462 XA8.XA4.MN0.G a_21080_45508# 6.57e-19
C9463 XA6.XA6.MP0.G XA6.XA1.XA2.MP0.D 0.0126f
C9464 XA3.XA1.XA5.MN2.G a_7328_42340# 1.97e-19
C9465 a_21080_46916# XA8.XA3.MN0.G 0.0658f
C9466 XA2.XA3.MN0.G XA3.XA3.MN0.G 1.48f
C9467 a_9848_46916# a_9848_46564# 0.0109f
C9468 D<1> XA7.XA1.XA4.MN1.D 0.00188f
C9469 XA3.XA4.MN0.D EN 0.0617f
C9470 VREF XA1.XA1.XA5.MP1.D 0.00623f
C9471 CK_SAMPLE a_21080_51140# 0.00759f
C9472 XA7.XA10.MP0.G a_18560_52548# 0.13f
C9473 AVDD a_2288_50788# 0.363f
C9474 SAR_IN XB1.M1.G 4.38e-19
C9475 XB2.XA1.MP0.D a_14960_2446# 0.00356f
C9476 a_14960_2798# XB2.XA4.MP0.D 0.00553f
C9477 XA20.XA3a.MN0.D a_13520_43044# 0.0905f
C9478 SARN li_14804_31260# 0.00103f
C9479 XA5.XA6.MP0.G XA5.XA1.XA1.MN0.D 0.00112f
C9480 D<5> a_7328_39876# 7.77e-20
C9481 a_11000_45156# a_12368_45156# 8.89e-19
C9482 XA2.XA1.XA5.MN2.D a_5960_44804# 0.156f
C9483 D<1> a_17408_40228# 3.45e-20
C9484 XA8.XA9.MN1.G a_19928_50788# 0.015f
C9485 AVDD a_4808_47972# 0.00125f
C9486 XA3.XA9.MN1.G a_7328_50436# 7.76e-19
C9487 XA5.XA7.MP0.D D<3> 2.65e-19
C9488 a_5960_51844# D<6> 1.25e-19
C9489 a_9848_51492# XA5.XA1.XA5.MN2.G 0.0674f
C9490 XDAC2.XC64b<1>.XRES1A.B XDAC2.X16ab.XRES1B.B 0.617f
C9491 a_17408_43748# a_18560_43748# 0.00133f
C9492 XA0.XA1.XA5.MN1.D a_n232_43396# 0.00176f
C9493 EN a_920_43396# 0.162f
C9494 XA20.XA3a.MN0.D a_12368_40580# 0.0658f
C9495 XA20.XA2a.MN0.D a_19928_41636# 0.0147f
C9496 AVDD a_18560_44804# 0.00125f
C9497 D<6> XA1.XA4.MN0.D 6.18f
C9498 XA0.XA6.MP0.G XA4.XA6.MP0.G 0.0763f
C9499 a_920_50436# a_920_50084# 0.0109f
C9500 XA1.XA6.MP0.G XA3.XA6.MP0.G 0.0635f
C9501 XA3.XA1.XA5.MN2.G a_5960_49028# 0.00363f
C9502 XDAC1.XC64a<0>.XRES8.B li_9184_10992# 9.91e-20
C9503 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES2.B 0.0307f
C9504 li_14804_11604# li_14804_10992# 0.00271f
C9505 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES16.B 0.0381f
C9506 XA2.XA1.XA4.MP1.D a_5960_42340# 0.00176f
C9507 a_18560_42692# a_19928_42692# 8.89e-19
C9508 EN a_n232_40932# 0.00712f
C9509 XA7.XA1.XA5.MN2.G a_16040_45860# 0.00363f
C9510 D<6> a_4808_46212# 0.0141f
C9511 a_920_49028# a_920_48676# 0.0109f
C9512 AVDD a_3440_42340# 0.00125f
C9513 D<2> a_16040_46564# 0.0695f
C9514 AVDD XA0.XA12.MP0.D 1.89f
C9515 a_17408_54308# a_18560_54308# 0.00133f
C9516 a_4808_54308# a_4808_53956# 0.0109f
C9517 a_4808_41284# a_5960_41284# 0.00133f
C9518 SARP li_9184_20820# 0.00103f
C9519 AVDD a_14960_2798# 0.465f
C9520 D<3> XA5.XA1.XA5.MN0.D 0.00188f
C9521 XA5.XA4.MN0.G a_12368_46564# 3.46e-19
C9522 a_21080_47620# a_21080_47268# 0.0109f
C9523 D<7> a_2288_43396# 7.77e-20
C9524 VREF a_17408_45156# 0.0195f
C9525 XA8.XA11.MN1.G XA8.XA9.MN1.G 0.00804f
C9526 XA3.XA11.MN1.G a_8480_52196# 5.56e-19
C9527 a_n232_52900# a_920_52900# 0.00133f
C9528 AVDD a_8480_51492# 0.00166f
C9529 CK_SAMPLE a_3440_51844# 2.08e-19
C9530 a_14888_39876# a_16040_39876# 0.00133f
C9531 XA5.XA1.XA5.MN2.G a_11000_40580# 0.0506f
C9532 XA2.XA3.MN0.G a_3440_44452# 2.51e-19
C9533 XA1.XA3.MN0.G a_4808_44452# 4.4e-20
C9534 XA4.XA4.MN0.G XA4.XA1.XA2.MP0.D 0.206f
C9535 XA0.XA4.MN0.D XA0.XA1.XA4.MP0.D 7.95e-19
C9536 XA20.XA3a.MN0.D a_8480_43748# 0.00228f
C9537 a_16040_45860# a_16040_45508# 0.0109f
C9538 XA20.XA2a.MN0.D a_22448_45156# 0.00407f
C9539 a_9848_51844# a_11000_51844# 0.00133f
C9540 XA3.XA7.MP0.D XA3.XA8.MP0.D 0.124f
C9541 XA6.XA9.MN1.G XA6.XA1.XA5.MN2.G 4.35e-19
C9542 AVDD a_2288_49028# 0.356f
C9543 CK_SAMPLE XA0.XA4.MN0.D 0.0364f
C9544 XA2.XA9.MN1.G a_4808_51140# 0.0469f
C9545 SARN a_23600_51492# 0.157f
C9546 a_19928_44100# EN 0.00576f
C9547 XA7.XA1.XA5.MN2.D a_17408_43396# 4.58e-19
C9548 XA20.XA2a.MN0.D XA2.XA1.XA4.MN0.D 0.0375f
C9549 XA0.XA1.XA5.MN2.D a_920_43044# 1.88e-19
C9550 D<7> li_9184_26556# 0.00504f
C9551 D<7> XA1.XA6.MN0.D 0.00148f
C9552 AVDD a_17408_45860# 0.356f
C9553 a_12368_50788# a_13520_50788# 0.00133f
C9554 XA5.XA6.MN2.D a_13520_50436# 0.00176f
C9555 XA3.XA1.XA5.MN2.G a_5960_50084# 0.00366f
C9556 a_16040_51844# VREF 0.00396f
C9557 a_9848_43044# XA4.XA1.XA4.MN1.D 0.00176f
C9558 XA1.XA1.XA2.MP0.D a_3440_42340# 0.0966f
C9559 XA5.XA1.XA2.MP0.D XA5.XA1.XA4.MP0.D 4.34e-19
C9560 EN a_5960_41636# 0.00649f
C9561 AVDD a_11000_43044# 0.381f
C9562 XA4.XA4.MN0.D XA5.XA4.MN0.D 0.00869f
C9563 XA0.XA4.MN0.D a_920_49380# 0.154f
C9564 VREF a_n232_49380# 8.08e-19
C9565 a_21080_41988# a_21080_41636# 0.0109f
C9566 XA6.XA6.MP0.G XA6.XA1.XA5.MN2.D 0.0325f
C9567 XA3.XA6.MP0.G a_7328_45156# 5.5e-19
C9568 XA4.XA1.XA5.MN2.G a_8480_43748# 2.66e-19
C9569 XA3.XA1.XA5.MN2.G a_9848_43748# 7.1e-20
C9570 XA4.XA4.MN0.G a_11000_47620# 0.155f
C9571 XA4.XA4.MN0.D a_9848_46212# 1.1e-19
C9572 VREF a_14888_46212# 7.12e-19
C9573 AVDD a_9848_40580# 0.00125f
C9574 a_14888_47972# a_16040_47972# 0.00133f
C9575 XA0.XA6.MP2.G EN 0.0666f
C9576 D<4> a_9848_44100# 6.49e-19
C9577 a_2288_47972# a_2288_47620# 0.0109f
C9578 AVDD XA6.XA9.MN1.G 0.93f
C9579 XA2.XA12.MP0.G a_4808_52900# 0.00258f
C9580 XA3.XA11.MN1.G a_5960_52900# 0.00183f
C9581 a_n232_53604# XA0.XA10.MP0.D 1.17e-19
C9582 a_12368_53604# a_12368_53252# 0.0109f
C9583 XA0.XA11.MN1.G a_n232_53252# 0.0689f
C9584 XA7.XA11.MN1.G XA7.XA10.MP0.D 0.0909f
C9585 XA6.XA12.MP0.G XA6.XA10.MP0.D 0.0632f
C9586 a_8480_40580# a_8480_40228# 0.0109f
C9587 XA0.XA6.MP0.G XA0.XA1.XA4.MP0.D 9.97e-19
C9588 a_8480_46212# a_9848_46212# 8.89e-19
C9589 a_22448_46564# a_22448_46212# 0.0109f
C9590 XA8.XA3.MN0.G a_21080_45860# 0.155f
C9591 XA1.XA3.MN0.G a_4808_45508# 4.4e-20
C9592 XA2.XA3.MN0.G a_3440_45508# 4.21e-19
C9593 XA7.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S 0.327f
C9594 XA0.XA7.MP0.G a_n232_41284# 0.00527f
C9595 XA4.XA6.MP0.G a_11000_42692# 5.5e-19
C9596 XA2.XA4.MN0.D a_5960_43396# 9.14e-20
C9597 XA1.XA4.MN0.G a_3440_44100# 0.0164f
C9598 XA8.XA4.MN0.G a_19928_44452# 0.00907f
C9599 XA6.XA9.MN1.G a_13520_52196# 2.84e-19
C9600 CK_SAMPLE XA0.XA6.MP0.G 0.046f
C9601 XA8.XA10.MP0.G a_19928_51844# 5.59e-19
C9602 XA2.XA10.MP0.G XA2.XA8.MP0.D 0.0434f
C9603 XA1.XA9.MN1.G XA1.XA7.MP0.D 0.274f
C9604 AVDD a_2288_50084# 0.358f
C9605 XB1.XA0.MP0.D a_9560_n18# 6.02e-19
C9606 XB1.XA3.MN0.S CK_SAMPLE_BSSW 0.00496f
C9607 XB2.XA3.MN0.S a_13808_686# 0.0328f
C9608 a_13808_1390# a_13808_1038# 0.0109f
C9609 XA4.XA4.MN0.G a_11000_41988# 5.1e-20
C9610 XA3.XA6.MP0.G a_11000_39876# 3.21e-19
C9611 a_16040_44804# a_16040_44452# 0.0109f
C9612 a_8480_45156# EN 4.58e-19
C9613 XA2.XA4.MN0.D a_4808_40932# 9.25e-20
C9614 SARN XDAC2.XC128b<2>.XRES2.B 6.99f
C9615 XA20.XA3a.MN0.D a_4808_42340# 0.00547f
C9616 XA5.XA1.XA5.MN2.D XA5.XA1.XA5.MP1.D 0.0488f
C9617 XA20.XA2a.MN0.D a_13520_43396# 4.8e-20
C9618 a_2288_44452# a_3440_44452# 0.00133f
C9619 XA3.XA1.XA5.MN2.G a_4808_50788# 1.87e-19
C9620 XA8.XA7.MP0.G XA8.XA6.MN2.D 6.33e-19
C9621 a_12368_52548# VREF 0.00396f
C9622 AVDD a_16040_46916# 0.359f
C9623 XA8.XA9.MN1.G a_19928_50084# 0.00969f
C9624 XB1.XA3.MN1.D m3_n2104_3300# 0.17f
C9625 XB2.XA4.MP0.D m3_25976_4356# 0.0137f
C9626 XDAC1.XC128b<2>.XRES8.B XDAC1.XC128b<2>.XRES2.B 0.44f
C9627 XDAC2.XC128b<2>.XRES8.B li_14804_21432# 9.91e-20
C9628 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES16.B 0.0483f
C9629 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES1A.B 0.00438f
C9630 XA0.XA6.MP0.G li_14804_15696# 1.85e-20
C9631 XA20.XA2a.MN0.D a_12368_40932# 0.0662f
C9632 XA6.XA1.XA5.MP0.D a_14888_43396# 2.16e-19
C9633 XA6.XA1.XA5.MN0.D a_16040_43396# 2.16e-19
C9634 a_2288_43396# a_3440_43396# 0.00133f
C9635 EN a_16040_42692# 0.159f
C9636 XA0.XA6.MP0.G a_920_49380# 0.0781f
C9637 XA4.XA1.XA5.MN2.G a_5960_47972# 7.1e-20
C9638 XA3.XA1.XA5.MN2.G a_7328_47972# 7.1e-20
C9639 AVDD a_5960_43748# 0.357f
C9640 XA3.XA6.MP0.D VREF 0.0115f
C9641 XA3.XA6.MP0.G XA1.XA4.MN0.D 1.9e-19
C9642 XA6.XA6.MN0.D a_14888_49732# 0.00176f
C9643 XA6.XA6.MP0.G a_16040_49732# 0.101f
C9644 li_9184_6288# li_9184_5676# 0.00271f
C9645 XA6.XA1.XA2.MP0.D a_16040_40932# 4.25e-20
C9646 XA5.XA1.XA4.MN0.D a_13520_41988# 0.00176f
C9647 a_13520_42340# a_14888_42340# 8.89e-19
C9648 VREF a_13520_47268# 1.19e-19
C9649 XA4.XA4.MN0.D a_8480_47268# 4.76e-20
C9650 XA3.XA4.MN0.D a_9848_47268# 4.76e-20
C9651 AVDD XA6.XA1.XA1.MP2.D 0.127f
C9652 D<3> XA5.XA1.XA5.MN2.D 0.0348f
C9653 D<0> a_19928_45508# 0.00245f
C9654 a_19928_48676# a_19928_48324# 0.0109f
C9655 a_9848_48676# XA4.XA4.MN0.G 1.34e-19
C9656 D<6> a_5960_45156# 6.68e-19
C9657 XA7.XA1.XA5.MN2.G a_16040_44804# 0.00486f
C9658 XA20.XA9.MP0.D a_23600_43044# 0.0714f
C9659 a_11000_53956# a_11000_53604# 0.0109f
C9660 CK_SAMPLE a_23600_53604# 7.07e-19
C9661 XA5.XA11.MN1.G XA4.XA12.MP0.G 0.142f
C9662 AVDD XA1.XA10.MP0.D 0.727f
C9663 a_23600_53956# XA20.XA10.MN0.D 0.00176f
C9664 XA0.XA1.XA1.MN0.D a_920_40580# 8.3e-19
C9665 XA5.XA1.XA1.MN0.D a_12368_40932# 8.29e-20
C9666 a_920_40932# a_2288_40932# 8.89e-19
C9667 SARP XDAC1.XC64a<0>.XRES2.B 6.99f
C9668 XA8.XA4.MN0.G a_19928_45508# 0.0104f
C9669 XA2.XA4.MN0.G XA2.XA1.XA5.MN2.D 0.135f
C9670 D<1> XA7.XA1.XA4.MP1.D 7.43e-19
C9671 XA3.XA1.XA5.MN2.G a_5960_42340# 0.00442f
C9672 a_19928_46916# XA8.XA3.MN0.G 0.0682f
C9673 XA1.XA3.MN0.G XA3.XA3.MN0.G 0.171f
C9674 XA2.XA4.MN0.D EN 0.0618f
C9675 VREF XA0.XA1.XA5.MP1.D 0.00623f
C9676 AVDD a_920_50788# 0.363f
C9677 CK_SAMPLE a_19928_51140# 0.0772f
C9678 a_5960_52548# a_7328_52548# 8.89e-19
C9679 XA7.XA10.MP0.G a_17408_52548# 0.0684f
C9680 XA0.XA10.MP0.G XA0.XA9.MN0.D 0.106f
C9681 a_13520_52900# XA5.XA9.MN1.G 0.00113f
C9682 XB2.XA1.MP0.D a_13808_2446# 0.0914f
C9683 a_9560_2446# a_11000_2446# 8e-19
C9684 SAR_IP XB1.XA4.MP0.D 0.00603f
C9685 a_8408_3502# XB1.XA3.MN1.D 1.93e-19
C9686 XA20.XA3a.MN0.D a_12368_43044# 0.00877f
C9687 XA2.XA1.XA5.MN2.D a_4808_44804# 0.153f
C9688 XA6.XA4.MN0.G XA6.XA1.XA4.MP1.D 0.0488f
C9689 XA0.XA4.MN0.G a_920_42692# 0.00224f
C9690 XA5.XA3.MN0.G a_13520_43748# 2.78e-19
C9691 AVDD a_3440_47972# 0.00125f
C9692 a_920_51492# a_920_51140# 0.0109f
C9693 a_18560_51492# a_19928_51492# 8.89e-19
C9694 XA8.XA11.MP0.D VREF 0.00246f
C9695 EN a_n232_43396# 0.00742f
C9696 XA2.XA3.MN0.G a_4808_41284# 0.00335f
C9697 XA20.XA3a.MN0.D a_11000_40580# 0.0674f
C9698 XA20.XA2a.MN0.D a_18560_41636# 0.0145f
C9699 XA5.XA1.XA5.MN1.D XA5.XA1.XA2.MP0.D 0.0102f
C9700 XA5.XA1.XA5.MP1.D XA5.XA1.XA5.MP0.D 0.0488f
C9701 a_3440_43748# XA1.XA1.XA5.MN0.D 0.00176f
C9702 AVDD a_17408_44804# 0.356f
C9703 a_16040_50436# XA6.XA6.MP0.G 0.0662f
C9704 a_14888_50436# XA6.XA6.MN0.D 0.00176f
C9705 D<6> VREF 1.3f
C9706 D<7> XA3.XA4.MN0.D 0.00195f
C9707 XA8.XA7.MP0.G a_22448_49380# 8.22e-19
C9708 XA7.XA1.XA4.MP1.D XA7.XA1.XA4.MP0.D 0.0488f
C9709 XA7.XA1.XA2.MP0.D a_18560_41636# 0.00316f
C9710 a_5960_42692# XA2.XA1.XA4.MP0.D 0.00176f
C9711 D<8> XDAC2.XC0.XRES2.B 0.00406f
C9712 a_12368_49028# a_13520_49028# 0.00133f
C9713 AVDD a_2288_42340# 0.361f
C9714 VREF a_12368_48324# 0.0536f
C9715 XA3.XA4.MN0.D a_8480_48324# 0.0997f
C9716 D<2> a_14888_46564# 0.0551f
C9717 AVDD a_23600_53956# 0.00159f
C9718 XA6.XA1.XA1.MP2.D a_16040_41284# 0.0465f
C9719 AVDD a_13808_2798# 0.00165f
C9720 D<3> XA5.XA1.XA5.MP0.D 7.43e-19
C9721 a_7328_47268# a_8480_47268# 0.00133f
C9722 XA5.XA1.XA5.MN2.G a_11000_43044# 0.00551f
C9723 XA1.XA6.MP0.G EN 0.065f
C9724 VREF a_16040_45156# 0.0195f
C9725 XA3.XA11.MN1.G a_7328_52196# 7.34e-19
C9726 a_18560_53252# a_18560_52900# 0.0109f
C9727 XA3.XA10.MP0.D a_8480_52900# 0.13f
C9728 XA8.XA11.MN1.G XA7.XA9.MN0.D 1.71e-19
C9729 AVDD a_7328_51492# 0.387f
C9730 XA8.XA3.MN0.G a_21080_44804# 0.00498f
C9731 XA1.XA3.MN0.G a_3440_44452# 0.0963f
C9732 XA4.XA1.XA5.MN2.G a_11000_40580# 5.68e-19
C9733 XA5.XA1.XA5.MN2.G a_9848_40580# 9.75e-19
C9734 SARN a_13808_2446# 0.00101f
C9735 XA0.XA4.MN0.D XA0.XA1.XA4.MN0.D 8.13e-19
C9736 XA20.XA3a.MN0.D a_7328_43748# 0.00106f
C9737 a_2288_45508# a_3440_45508# 0.00133f
C9738 AVDD a_920_49028# 0.356f
C9739 XA8.XA7.MP0.D a_21080_51844# 0.133f
C9740 a_22448_54308# VREF 0.0013f
C9741 XA2.XA9.MN1.G a_3440_51140# 2.84e-19
C9742 XA5.XA9.MN1.G XA7.XA1.XA5.MN2.G 4.35e-19
C9743 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES1A.B 0.00438f
C9744 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES16.B 0.0483f
C9745 XDAC2.XC0.XRES8.B XDAC2.XC0.XRES2.B 0.44f
C9746 SARN li_14804_10992# 0.00103f
C9747 XA20.XA3a.MN0.D XA7.XA1.XA1.MN0.S 0.0673f
C9748 a_18560_44100# EN 0.00576f
C9749 a_21080_44100# a_22448_44100# 8.89e-19
C9750 XA20.XA2a.MN0.D XA1.XA1.XA4.MN0.D 0.0409f
C9751 XA0.XA1.XA5.MN2.D a_n232_43044# 5.1e-20
C9752 XA0.XA6.MP2.G XDAC1.X16ab.XRES1B.B 4.06e-21
C9753 a_8480_44100# XA3.XA1.XA5.MN1.D 0.00176f
C9754 XA8.XA7.MP0.G XA20.XA3.MN6.D 0.256f
C9755 D<7> XA1.XA6.MP0.D 0.0323f
C9756 AVDD a_16040_45860# 0.356f
C9757 a_n232_50788# a_n232_50436# 0.0109f
C9758 XDAC2.XC128a<1>.XRES8.B XDAC2.XC32a<0>.XRES8.B 6.7e-19
C9759 li_14804_16728# li_14804_16116# 0.00271f
C9760 EN a_4808_41636# 1.25e-19
C9761 XA0.XA4.MN0.D li_9184_15696# 1.85e-20
C9762 XA1.XA1.XA2.MP0.D a_2288_42340# 2.54e-19
C9763 a_21080_43044# a_22448_43044# 8.89e-19
C9764 a_12368_49732# a_12368_49380# 0.0109f
C9765 XA2.XA6.MP0.G a_5960_48324# 0.00417f
C9766 VREF XA8.XA4.MN0.D 0.588f
C9767 XA0.XA4.MN0.D a_n232_49380# 0.155f
C9768 XA6.XA6.MP0.G a_16040_48676# 0.0881f
C9769 AVDD a_9848_43044# 0.00125f
C9770 a_21080_42340# XA8.XA1.XA1.MN0.S 1.34e-19
C9771 a_7328_41636# a_8480_41636# 0.00133f
C9772 SARP li_9184_31260# 0.00103f
C9773 XA3.XA1.XA5.MN2.G a_8480_43748# 0.0749f
C9774 XA4.XA1.XA5.MN2.G a_7328_43748# 0.00442f
C9775 XA4.XA4.MN0.G a_9848_47620# 0.154f
C9776 VREF a_13520_46212# 7.12e-19
C9777 AVDD a_8480_40580# 0.00125f
C9778 AVDD XA5.XA9.MN0.D 4.25e-19
C9779 CK_SAMPLE XA20.XA4.MN0.D 0.0115f
C9780 XA7.XA11.MN1.G XA6.XA10.MP0.D 0.00744f
C9781 a_19928_40580# a_21080_40580# 0.00133f
C9782 XA20.XA3a.MN0.D a_18560_44804# 1.57e-20
C9783 SARN a_23600_40580# 8.72e-19
C9784 XA0.XA6.MP0.G XA0.XA1.XA4.MN0.D 6.07e-19
C9785 XA1.XA3.MN0.G a_3440_45508# 0.109f
C9786 XA8.XA3.MN0.G a_19928_45860# 0.162f
C9787 XA6.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S 0.0308f
C9788 XA4.XA6.MP0.G a_9848_42692# 7.76e-20
C9789 XA2.XA4.MN0.D a_4808_43396# 9.25e-20
C9790 VREF a_7328_43396# 3.39e-19
C9791 XA1.XA4.MN0.G a_2288_44100# 6.11e-19
C9792 XA7.XA4.MN0.G a_19928_44452# 2.2e-19
C9793 XA8.XA4.MN0.G a_18560_44452# 2.2e-19
C9794 a_920_52196# a_2288_52196# 8.89e-19
C9795 a_18560_52548# XA7.XA7.MP0.D 5.16e-20
C9796 XA5.XA9.MN0.D a_13520_52196# 0.0492f
C9797 XA5.XA9.MN1.G a_14888_52196# 2.84e-19
C9798 AVDD a_920_50084# 0.358f
C9799 XB2.XA0.MP0.D a_14960_334# 0.00524f
C9800 XB1.XA0.MP0.D a_8408_n18# 0.00102f
C9801 a_8408_1038# a_9560_1038# 0.00133f
C9802 XA4.XA4.MN0.G a_9848_41988# 1.74e-19
C9803 XA3.XA6.MP0.G a_9848_39876# 8.95e-19
C9804 a_7328_45156# EN 1.83e-19
C9805 XA20.XA3a.MN0.D a_3440_42340# 0.00552f
C9806 a_11000_51140# XA4.XA6.MP2.D 0.00176f
C9807 XA0.XA6.MP2.G D<7> 2.22f
C9808 a_11000_52548# VREF 0.00396f
C9809 AVDD a_14888_46916# 0.00131f
C9810 XA8.XA7.MP0.G D<0> 0.6f
C9811 XB2.XA4.MP0.D m3_16544_4532# 0.0634f
C9812 XB1.XA3.MN1.D m3_7544_3476# 0.0137f
C9813 XA20.XA2a.MN0.D a_11000_40932# 0.0678f
C9814 XA2.XA1.XA2.MP0.D a_5960_43044# 3.59e-19
C9815 XA2.XA1.XA5.MN0.D a_4808_43044# 0.00176f
C9816 XA6.XA1.XA5.MN0.D a_14888_43396# 0.0474f
C9817 XA0.XA6.MP0.G a_n232_49380# 0.0547f
C9818 XA3.XA1.XA5.MN2.G a_5960_47972# 0.00363f
C9819 XA2.XA6.MP0.G XA3.XA4.MN0.D 0.0657f
C9820 XA8.XA7.MP0.G XA8.XA4.MN0.G 0.158f
C9821 AVDD a_4808_43748# 0.00125f
C9822 XA3.XA6.MP0.G VREF 0.568f
C9823 XA6.XA6.MP0.G a_14888_49732# 0.00239f
C9824 a_n232_50084# a_n232_49732# 0.0109f
C9825 a_12368_50084# a_13520_50084# 0.00133f
C9826 SARP a_13808_2446# 2.97e-20
C9827 D<8> li_14804_21432# 3.5e-20
C9828 a_920_42692# XA0.XA1.XA1.MN0.S 6.76e-20
C9829 a_920_42340# a_920_41988# 0.0109f
C9830 XA3.XA4.MN0.D a_8480_47268# 0.0963f
C9831 VREF a_12368_47268# 0.0191f
C9832 a_5960_48324# a_7328_48324# 8.89e-19
C9833 D<6> a_4808_45156# 7.77e-19
C9834 XA7.XA1.XA5.MN2.G a_14888_44804# 1.86e-19
C9835 XA20.XA9.MP0.D a_22448_43044# 0.139f
C9836 AVDD XA6.XA1.XA1.MN0.S 1.04f
C9837 XA3.XA12.MP0.G XA4.XA12.MP0.G 0.00217f
C9838 CK_SAMPLE a_22448_53604# 0.00904f
C9839 XA4.XA11.MN1.G XA6.XA11.MN1.G 1.54e-19
C9840 AVDD XA0.XA10.MP0.D 0.728f
C9841 a_23600_53956# XA20.XA10.MN1.D 0.0314f
C9842 XA0.XA1.XA1.MN0.D a_n232_40580# 0.035f
C9843 XA5.XA1.XA1.MP1.D a_12368_40932# 0.0465f
C9844 a_8480_46916# a_8480_46564# 0.0109f
C9845 XA8.XA4.MN0.G a_18560_45508# 2.84e-19
C9846 XA7.XA4.MN0.G a_19928_45508# 2.84e-19
C9847 XA2.XA4.MN0.G XA1.XA1.XA5.MN2.D 0.0024f
C9848 XA1.XA4.MN0.G XA2.XA1.XA5.MN2.D 0.0024f
C9849 XA3.XA1.XA5.MN2.G a_4808_42340# 3.12e-19
C9850 XA1.XA3.MN0.G XA2.XA3.MN0.G 3.47f
C9851 D<8> XA3.XA3.MN0.G 0.216f
C9852 XA8.XA7.MP0.G XA8.XA1.XA4.MP0.D 0.00358f
C9853 XA2.XA1.XA5.MN2.G a_5960_42340# 1.97e-19
C9854 D<5> a_8480_42692# 6.49e-19
C9855 XA0.XA4.MN0.D XA0.XA1.XA5.MP1.D 9.69e-19
C9856 XA1.XA4.MN0.D EN 0.0617f
C9857 AVDD a_n232_50788# 0.00154f
C9858 CK_SAMPLE a_18560_51140# 0.067f
C9859 XA0.XA10.MP0.G XA0.XA9.MN1.G 0.202f
C9860 a_14960_2798# XB2.M1.G 4.74e-19
C9861 SAR_IP XB1.M1.G 0.679f
C9862 XB2.XA1.MN0.D a_14960_2446# 0.0674f
C9863 XB1.XA1.MN0.D XB1.XA4.MP0.D 0.0122f
C9864 XB1.XA1.MP0.D XB1.XA4.MN0.D 0.0109f
C9865 XB2.XA1.MP0.D a_12368_2446# 3.77e-19
C9866 SAR_IN a_13808_2446# 1.82e-19
C9867 XA20.XA3a.MN0.D a_11000_43044# 0.00835f
C9868 SARN XDAC2.XC0.XRES2.B 6.99f
C9869 a_9848_45156# a_11000_45156# 0.00133f
C9870 XA1.XA6.MP0.G a_3440_40932# 3.97e-20
C9871 XA6.XA4.MN0.G XA6.XA1.XA4.MN1.D 0.0642f
C9872 XA0.XA4.MN0.G a_n232_42692# 0.0049f
C9873 XA3.XA4.MN0.D a_8480_41636# 9.24e-20
C9874 AVDD a_2288_47972# 0.356f
C9875 a_8480_51492# XA4.XA1.XA5.MN2.G 0.0658f
C9876 XA7.XA11.MP0.D VREF 0.00176f
C9877 XDAC1.XC64b<1>.XRES1A.B XDAC1.X16ab.XRES1B.B 0.617f
C9878 XA2.XA3.MN0.G a_3440_41284# 4.21e-19
C9879 XA1.XA3.MN0.G a_4808_41284# 4.4e-20
C9880 EN XA8.XA1.XA5.MP0.D 0.0426f
C9881 D<6> XDAC1.XC128a<1>.XRES16.B 3.2e-20
C9882 XA0.XA6.MP2.G li_9184_16116# 0.00508f
C9883 XA20.XA3a.MN0.D a_9848_40580# 0.0658f
C9884 XA20.XA2a.MN0.D a_17408_41636# 0.00184f
C9885 XA5.XA1.XA5.MP1.D XA5.XA1.XA2.MP0.D 6.52e-20
C9886 a_16040_43748# a_17408_43748# 8.89e-19
C9887 a_n232_50436# a_n232_50084# 0.0109f
C9888 a_14888_50436# XA6.XA6.MP0.G 3.02e-20
C9889 D<7> XA2.XA4.MN0.D 0.00522f
C9890 D<6> XA0.XA4.MN0.D 0.293f
C9891 XA8.XA7.MP0.G a_21080_49380# 0.00363f
C9892 D<3> a_13520_49732# 7.01e-19
C9893 AVDD a_16040_44804# 0.356f
C9894 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES2.B 0.0307f
C9895 li_9184_11604# li_9184_10992# 0.00271f
C9896 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES16.B 0.0381f
C9897 SARP a_23600_40580# 0.0717f
C9898 XA3.XA1.XA2.MP0.D XA3.XA1.XA1.MN0.S 2.11e-19
C9899 XA7.XA1.XA2.MP0.D a_17408_41636# 0.00224f
C9900 XA2.XA1.XA4.MN1.D a_4808_42340# 0.00176f
C9901 a_17408_42692# a_18560_42692# 0.00133f
C9902 D<8> XDAC1.XC0.XRES2.B 1.94e-19
C9903 a_n232_49028# a_n232_48676# 0.0109f
C9904 XA6.XA6.MP0.G a_16040_47620# 6.35e-19
C9905 AVDD a_920_42340# 0.361f
C9906 VREF a_11000_48324# 0.0536f
C9907 XA3.XA4.MN0.D a_7328_48324# 0.0682f
C9908 D<5> XA20.XA2a.MN0.D 0.076f
C9909 XA2.XA6.MP0.G a_5960_47268# 5.95e-19
C9910 AVDD a_22448_53956# 0.405f
C9911 a_16040_54308# a_17408_54308# 8.89e-19
C9912 a_3440_54308# a_3440_53956# 0.0109f
C9913 SARP XDAC1.XC128b<2>.XRES2.B 6.99f
C9914 XA1.XA1.XA1.MP2.D XA1.XA1.XA1.MP1.D 0.0488f
C9915 XA1.XA1.XA1.MN0.S XA1.XA1.XA1.MN0.D 0.0743f
C9916 a_3440_41284# a_4808_41284# 8.89e-19
C9917 XA6.XA1.XA1.MN0.S a_16040_41284# 0.0964f
C9918 D<3> XA5.XA1.XA2.MP0.D 0.0153f
C9919 XA0.XA6.MP0.G XA0.XA1.XA5.MP1.D 0.00121f
C9920 XA4.XA4.MN0.G a_11000_46564# 3.46e-19
C9921 a_19928_47620# a_19928_47268# 0.0109f
C9922 XA5.XA1.XA5.MN2.G a_9848_43044# 2.31e-19
C9923 VREF a_14888_45156# 7.39e-19
C9924 XA3.XA11.MN1.G a_5960_52196# 4.29e-19
C9925 XA3.XA10.MP0.D a_7328_52900# 0.0877f
C9926 XA8.XA11.MN1.G XA7.XA9.MN1.G 0.0169f
C9927 AVDD a_5960_51492# 0.387f
C9928 a_13520_39876# a_14888_39876# 8.89e-19
C9929 XA8.XA3.MN0.G a_19928_44804# 0.0404f
C9930 XA1.XA3.MN0.G a_2288_44452# 0.055f
C9931 XA3.XA4.MN0.G XA3.XA1.XA5.MN0.D 0.0198f
C9932 XA6.XA6.MP0.G a_16040_41988# 5.5e-19
C9933 D<4> XA4.XA1.XA1.MN0.D 0.0192f
C9934 XA4.XA1.XA5.MN2.G a_9848_40580# 0.083f
C9935 SARN a_12368_2446# 0.0039f
C9936 XA2.XA6.MP0.G a_5960_41636# 5.5e-19
C9937 XA20.XA3a.MN0.D a_5960_43748# 0.00106f
C9938 a_14888_45860# a_14888_45508# 0.0109f
C9939 XA1.XA9.MN1.G a_4808_51140# 2.84e-19
C9940 AVDD a_n232_49028# 0.00154f
C9941 a_8480_51844# a_9848_51844# 8.89e-19
C9942 XA8.XA7.MP0.D a_19928_51844# 0.159f
C9943 XA2.XA7.MP0.D XA2.XA8.MP0.D 0.124f
C9944 a_21080_54308# VREF 0.00569f
C9945 CK_SAMPLE a_22448_49732# 3.39e-19
C9946 XA5.XA9.MN1.G XA6.XA1.XA5.MN2.G 0.0494f
C9947 a_17408_44100# EN 0.0767f
C9948 XA6.XA1.XA5.MN2.D a_16040_43396# 4.58e-19
C9949 XA20.XA2a.MN0.D XA1.XA1.XA4.MP0.D 0.0255f
C9950 a_8480_44804# XA3.XA1.XA2.MP0.D 2.6e-20
C9951 D<7> XDAC1.XC64b<1>.XRES1A.B 0.00405f
C9952 XA8.XA7.MP0.G XA20.XA3a.MN0.G 0.0152f
C9953 D<7> XA1.XA6.MP0.G 0.537f
C9954 AVDD a_14888_45860# 0.00125f
C9955 a_11000_50788# a_12368_50788# 8.89e-19
C9956 XA5.XA6.MP2.D a_12368_50436# 0.00176f
C9957 D<3> a_13520_50436# 5.7e-19
C9958 D<6> XA0.XA6.MP0.G 0.0695f
C9959 EN a_3440_41636# 1.25e-19
C9960 a_8480_43044# XA3.XA1.XA4.MN1.D 0.00176f
C9961 XA2.XA6.MP0.G a_4808_48324# 0.00295f
C9962 VREF XA7.XA4.MN0.D 0.593f
C9963 XA3.XA4.MN0.D XA4.XA4.MN0.D 0.00869f
C9964 XA6.XA6.MP0.G a_14888_48676# 0.0651f
C9965 AVDD a_8480_43044# 0.00125f
C9966 a_7328_41988# XA3.XA1.XA1.MN0.S 3.8e-19
C9967 a_19928_41988# a_19928_41636# 0.0109f
C9968 VREF a_12368_46212# 0.0671f
C9969 XA3.XA4.MN0.D a_8480_46212# 6.37e-19
C9970 AVDD a_7328_40580# 0.381f
C9971 a_13520_47972# a_14888_47972# 8.89e-19
C9972 SARN a_23600_43044# 0.00188f
C9973 a_920_47972# a_920_47620# 0.0109f
C9974 AVDD XA5.XA9.MN1.G 0.93f
C9975 XA20.XA10.MN0.D a_23600_53252# 0.00176f
C9976 CK_SAMPLE XA8.XA10.MP0.G 0.00465f
C9977 a_11000_53604# a_11000_53252# 0.0109f
C9978 a_7328_40580# a_7328_40228# 0.0109f
C9979 a_7328_46212# a_8480_46212# 0.00133f
C9980 a_21080_46564# a_21080_46212# 0.0109f
C9981 XA1.XA3.MN0.G a_2288_45508# 0.0682f
C9982 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MP2.D 0.0739f
C9983 XA5.XA1.XA5.MN2.G XA6.XA1.XA1.MN0.S 5.21e-19
C9984 XA0.XA11.MN1.G a_13808_1038# 0.00173f
C9985 VREF a_5960_43396# 3.39e-19
C9986 XA7.XA4.MN0.G a_18560_44452# 0.00907f
C9987 CK_SAMPLE a_22448_50436# 0.00141f
C9988 XA7.XA10.MP0.G a_18560_51844# 5.59e-19
C9989 XA0.XA9.MN0.D XA0.XA7.MP0.D 0.00986f
C9990 XA1.XA10.MP0.G XA1.XA8.MP0.D 0.0434f
C9991 XA5.XA9.MN1.G a_13520_52196# 0.0878f
C9992 AVDD a_n232_50084# 0.00144f
C9993 XB2.XA0.MP0.D a_13808_334# 0.00401f
C9994 a_12368_1390# a_12368_1038# 0.0109f
C9995 XA6.XA3.MN0.G a_14888_43044# 3.62e-20
C9996 XA3.XA6.MP0.G a_8480_39876# 9.73e-19
C9997 a_14888_44804# a_14888_44452# 0.0109f
C9998 a_5960_45156# EN 1.83e-19
C9999 XA7.XA6.MP0.G a_18560_40228# 3.45e-20
C10000 XA1.XA4.MN0.D a_3440_40932# 9.24e-20
C10001 SARN li_14804_21432# 0.00103f
C10002 XA4.XA1.XA5.MN2.D XA4.XA1.XA5.MP1.D 0.0488f
C10003 a_920_44452# a_2288_44452# 8.89e-19
C10004 AVDD a_13520_46916# 0.00131f
C10005 XA0.XA6.MP2.G XA0.XA6.MP2.D 0.0399f
C10006 XA2.XA1.XA5.MN2.G a_3440_50788# 1.87e-19
C10007 XA2.XA9.MN1.G a_5960_49732# 0.0215f
C10008 XB2.XA4.MP0.D m3_16472_4532# 0.106f
C10009 XB1.XA3.MN1.D m3_7472_3476# 0.0137f
C10010 li_14804_22044# li_14804_21432# 0.00271f
C10011 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES2.B 0.0307f
C10012 XDAC1.XC128b<2>.XRES8.B li_9184_21432# 9.91e-20
C10013 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES16.B 0.0381f
C10014 XDAC2.X16ab.XRES1A.B XDAC2.XC128b<2>.XRES1A.B 0.00444f
C10015 XA0.XA6.MP0.G XDAC2.XC32a<0>.XRES1B.B 2.23e-21
C10016 XA20.XA2a.MN0.D a_9848_40932# 0.0717f
C10017 XA2.XA1.XA2.MP0.D a_4808_43044# 0.0292f
C10018 a_920_43396# a_2288_43396# 8.89e-19
C10019 XA6.XA1.XA2.MP0.D a_14888_43396# 0.0945f
C10020 D<3> a_13520_48676# 3.48e-19
C10021 XA2.XA6.MP0.G XA2.XA4.MN0.D 4.49f
C10022 D<7> a_3440_48324# 6.53e-19
C10023 XA8.XA1.XA5.MN2.G XA8.XA4.MN0.G 0.168f
C10024 AVDD a_3440_43748# 0.00125f
C10025 XA2.XA6.MP0.D VREF 0.0115f
C10026 XA3.XA6.MP0.G XA0.XA4.MN0.D 1.36e-19
C10027 SARN XA3.XA3.MN0.G 0.0911f
C10028 XDAC2.XC1.XRES16.B XDAC2.XC1.XRES1A.B 0.454f
C10029 SARP a_12368_2446# 0.0418f
C10030 XA5.XA1.XA4.MP0.D a_12368_41988# 0.00176f
C10031 a_12368_42340# a_13520_42340# 0.00133f
C10032 XA3.XA4.MN0.D a_7328_47268# 0.0576f
C10033 VREF a_11000_47268# 0.0191f
C10034 XA2.XA6.MP0.G a_5960_46212# 5.5e-19
C10035 a_18560_48676# a_18560_48324# 0.0109f
C10036 a_8480_48676# XA3.XA4.MN0.G 1.34e-19
C10037 XA6.XA1.XA5.MN2.G a_14888_44804# 1.95e-19
C10038 XA20.XA9.MP0.D a_21080_43044# 5.7e-20
C10039 XA4.XA6.MP0.G XA20.XA2a.MN0.D 0.0783f
C10040 AVDD XA5.XA1.XA1.MP2.D 0.127f
C10041 XA4.XA11.MN1.G XA4.XA12.MP0.G 0.214f
C10042 a_9848_53956# a_9848_53604# 0.0109f
C10043 CK_SAMPLE a_21080_53604# 7.43e-19
C10044 AVDD a_23600_53252# 0.00166f
C10045 a_22448_53956# XA20.XA10.MN1.D 0.00224f
C10046 XA4.XA1.XA1.MN0.S a_11000_40228# 0.0313f
C10047 a_n232_40932# a_920_40932# 0.00133f
C10048 SARP li_9184_10992# 0.00103f
C10049 XA7.XA4.MN0.G a_18560_45508# 0.0104f
C10050 XA1.XA4.MN0.G XA1.XA1.XA5.MN2.D 0.135f
C10051 XA1.XA6.MP0.G a_3440_43396# 7.76e-20
C10052 XA8.XA1.XA5.MN2.G XA8.XA1.XA4.MP0.D 6.33e-19
C10053 a_18560_46916# XA7.XA3.MN0.G 0.0666f
C10054 D<8> XA2.XA3.MN0.G 0.0394f
C10055 XA8.XA7.MP0.G XA8.XA1.XA4.MN0.D 7.2e-19
C10056 XA2.XA1.XA5.MN2.G a_4808_42340# 0.00568f
C10057 D<5> a_7328_42692# 7.77e-20
C10058 XA0.XA4.MN0.D XA0.XA1.XA5.MN1.D 9.9e-19
C10059 VREF EN 0.911f
C10060 AVDD XA8.XA6.MP2.D 0.163f
C10061 CK_SAMPLE a_17408_51140# 8.45e-19
C10062 a_4808_52548# a_5960_52548# 0.00133f
C10063 XA6.XA10.MP0.G a_16040_52548# 0.07f
C10064 a_13808_2798# XB2.M1.G 0.00245f
C10065 a_8408_2446# a_9560_2446# 0.00133f
C10066 XB2.XA1.MN0.D a_13808_2446# 0.0711f
C10067 XB1.XA1.MN0.D XB1.M1.G 0.0319f
C10068 XB1.XA1.MP0.D XB1.XA4.MP0.D 0.0044f
C10069 a_8408_3854# XB1.XA3.MN1.D 1.93e-19
C10070 SAR_IN a_12368_2446# 0.0495f
C10071 XA20.XA3a.MN0.D a_9848_43044# 0.0864f
C10072 XA1.XA1.XA5.MN2.D a_3440_44804# 0.153f
C10073 XA8.XA1.XA5.MN2.D a_21080_45156# 0.155f
C10074 XA1.XA6.MP0.G a_2288_40932# 4.24e-19
C10075 XA3.XA4.MN0.D a_7328_41636# 9.15e-20
C10076 XA2.XA9.MN1.G a_5960_50436# 7.76e-19
C10077 AVDD a_920_47972# 0.356f
C10078 a_n232_51492# a_n232_51140# 0.0109f
C10079 a_7328_51492# XA4.XA1.XA5.MN2.G 0.0714f
C10080 XA7.XA9.MN1.G a_18560_50788# 0.015f
C10081 a_17408_51492# a_18560_51492# 0.00133f
C10082 XA6.XA11.MP0.D VREF 0.00185f
C10083 XA1.XA3.MN0.G a_3440_41284# 0.00342f
C10084 EN XA8.XA1.XA5.MN0.D 0.0044f
C10085 XA20.XA3a.MN0.D a_8480_40580# 0.0674f
C10086 XA20.XA2a.MN0.D a_16040_41636# 0.00184f
C10087 SARP a_23600_43044# 0.0855f
C10088 a_3440_43748# XA1.XA1.XA2.MP0.D 0.0686f
C10089 a_2288_43748# XA1.XA1.XA5.MP0.D 0.00176f
C10090 XA1.XA6.MP0.G XA2.XA6.MP0.G 2.62f
C10091 XA0.XA6.MP0.G XA3.XA6.MP0.G 0.0682f
C10092 XA1.XA6.MP2.D VREF 5.13e-19
C10093 D<7> XA1.XA4.MN0.D 6.79f
C10094 D<3> a_12368_49732# 0.0109f
C10095 AVDD a_14888_44804# 0.00125f
C10096 XA6.XA1.XA4.MP1.D XA6.XA1.XA4.MP0.D 0.0488f
C10097 a_4808_42692# XA2.XA1.XA4.MN0.D 0.00176f
C10098 D<8> li_14804_31872# 0.00508f
C10099 a_11000_49028# a_12368_49028# 8.89e-19
C10100 XA6.XA6.MP0.G a_14888_47620# 4.4e-19
C10101 AVDD a_n232_42340# 0.00125f
C10102 XA2.XA6.MP0.G a_4808_47268# 1.38e-19
C10103 AVDD a_21080_53956# 0.461f
C10104 XA1.XA1.XA1.MN0.S XA1.XA1.XA1.MP1.D 0.0615f
C10105 XA6.XA1.XA1.MN0.S a_14888_41284# 0.0658f
C10106 XA4.XA6.MP0.G a_11000_44100# 5.5e-19
C10107 XA0.XA6.MP0.G XA0.XA1.XA5.MN1.D 7.41e-19
C10108 XA4.XA4.MN0.G a_9848_46564# 0.0155f
C10109 a_5960_47268# a_7328_47268# 8.89e-19
C10110 XA4.XA1.XA5.MN2.G a_9848_43044# 0.0748f
C10111 VREF a_13520_45156# 7.39e-19
C10112 a_4808_53604# XA2.XA9.MN1.G 7.36e-20
C10113 XA7.XA11.MN1.G XA7.XA9.MN0.D 1.35e-19
C10114 a_17408_53252# a_17408_52900# 0.0109f
C10115 AVDD a_4808_51492# 0.00166f
C10116 CK_SAMPLE a_n232_51844# 1.64e-19
C10117 XA3.XA3.MN0.G SARP 0.0333f
C10118 XA3.XA4.MN0.G XA3.XA1.XA5.MP0.D 0.00138f
C10119 XA6.XA6.MP0.G a_14888_41988# 7.76e-20
C10120 XA4.XA1.XA5.MN2.G a_8480_40580# 0.00564f
C10121 XA3.XA1.XA5.MN2.G a_9848_40580# 7.1e-20
C10122 XA0.XA6.MP2.G a_920_40932# 4.07e-20
C10123 SARN a_11000_2446# 0.0438f
C10124 XA2.XA6.MP0.G a_4808_41636# 7.76e-20
C10125 XA20.XA3a.MN0.D a_4808_43748# 0.00218f
C10126 a_2288_45860# XA1.XA1.XA5.MN2.D 3.12e-20
C10127 a_920_45508# a_2288_45508# 8.89e-19
C10128 XA1.XA9.MN1.G a_3440_51140# 0.0469f
C10129 AVDD a_23600_49380# 0.00154f
C10130 CK_SAMPLE a_21080_49732# 5.27e-19
C10131 XDAC2.XC0.XRES8.B li_14804_31872# 9.91e-20
C10132 XDAC1.XC0.XRES8.B XDAC1.XC0.XRES2.B 0.44f
C10133 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES1A.B 0.00438f
C10134 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES16.B 0.0483f
C10135 a_16040_44100# EN 0.0752f
C10136 a_19928_44100# a_21080_44100# 0.00133f
C10137 SARN XDAC2.XC64a<0>.XRES8.B 27.7f
C10138 XA20.XA3a.MN0.D XA6.XA1.XA1.MN0.S 0.0673f
C10139 D<6> XDAC1.XC64b<1>.XRES16.B 3.2e-20
C10140 XA6.XA1.XA5.MN2.D a_14888_43396# 1.28e-19
C10141 XA20.XA2a.MN0.D XA0.XA1.XA4.MP0.D 0.0251f
C10142 a_18560_45156# XA7.XA1.XA2.MP0.D 1.56e-20
C10143 XA0.XA6.MP2.G li_9184_26556# 3.5e-20
C10144 XA3.XA3.MN0.G a_9848_42340# 7.54e-19
C10145 a_7328_44100# XA3.XA1.XA5.MP1.D 0.00176f
C10146 AVDD a_13520_45860# 0.00125f
C10147 D<3> a_12368_50436# 0.0863f
C10148 a_12368_51844# VREF 0.00396f
C10149 a_12368_51140# XA5.XA6.MP0.G 6.76e-20
C10150 li_9184_16728# li_9184_16116# 0.00271f
C10151 XDAC1.XC128a<1>.XRES8.B XDAC1.XC32a<0>.XRES8.B 6.7e-19
C10152 XA0.XA6.MP0.G li_14804_5676# 0.00506f
C10153 EN a_2288_41636# 0.00649f
C10154 XA0.XA4.MN0.D XDAC1.XC32a<0>.XRES1B.B 2.23e-21
C10155 a_19928_43044# a_21080_43044# 0.00133f
C10156 a_11000_49732# a_11000_49380# 0.0109f
C10157 XA20.XA3.MN0.D a_23600_49380# 0.0297f
C10158 VREF XA6.XA4.MN0.D 0.593f
C10159 D<3> a_13520_47620# 5.21e-19
C10160 D<7> a_3440_47268# 3.18e-19
C10161 XA6.XA1.XA5.MN2.G a_12368_46916# 0.00455f
C10162 AVDD a_7328_43044# 0.381f
C10163 a_5960_41636# a_7328_41636# 8.89e-19
C10164 SARP XDAC1.XC0.XRES2.B 6.99f
C10165 XA3.XA1.XA5.MN2.G a_5960_43748# 0.00442f
C10166 XA8.XA7.MP0.G XA8.XA1.XA5.MP1.D 0.00329f
C10167 XA3.XA4.MN0.G a_8480_47620# 0.154f
C10168 VREF a_11000_46212# 0.0671f
C10169 XA3.XA4.MN0.D a_7328_46212# 9.15e-20
C10170 AVDD a_5960_40580# 0.381f
C10171 AVDD XA4.XA9.MN0.D 4.25e-19
C10172 XA20.XA10.MN1.D a_23600_53252# 0.0865f
C10173 DONE a_23600_52548# 1.97e-19
C10174 XA1.XA12.MP0.G a_3440_52900# 0.00258f
C10175 XA2.XA11.MN1.G a_4808_52900# 7.39e-19
C10176 XA6.XA11.MN1.G XA6.XA10.MP0.D 0.0625f
C10177 XA5.XA12.MP0.G XA5.XA10.MP0.D 0.0632f
C10178 a_18560_40580# a_19928_40580# 8.89e-19
C10179 D<3> a_13520_41988# 6.49e-19
C10180 XA7.XA3.MN0.G a_18560_45860# 0.162f
C10181 D<7> a_3440_41636# 6.49e-19
C10182 XA6.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.S 0.301f
C10183 XA0.XA11.MN1.G a_12368_1038# 0.00151f
C10184 XA7.XA6.MP0.G XA7.XA1.XA4.MN1.D 7.41e-19
C10185 XA1.XA4.MN0.D a_3440_43396# 9.24e-20
C10186 XA0.XA4.MN0.G a_920_44100# 6.11e-19
C10187 XA7.XA4.MN0.G a_17408_44452# 5.54e-19
C10188 AVDD XA20.XA3.MN1.D 0.439f
C10189 CK_SAMPLE a_21080_50436# 0.00182f
C10190 a_n232_52196# a_920_52196# 0.00133f
C10191 XA0.XA9.MN1.G XA0.XA7.MP0.D 0.274f
C10192 XA5.XA9.MN1.G a_12368_52196# 0.0665f
C10193 XA7.XA10.MP0.G a_17408_51844# 0.00224f
C10194 XA3.XA4.MN0.G a_8480_41988# 1.74e-19
C10195 XA3.XA6.MP0.G a_7328_39876# 0.00207f
C10196 a_4808_45156# EN 4.58e-19
C10197 XA7.XA6.MP0.G a_17408_40228# 5.81e-19
C10198 XA1.XA4.MN0.D a_2288_40932# 9.15e-20
C10199 XA4.XA1.XA5.MN2.D XA4.XA1.XA5.MN1.D 0.0488f
C10200 XA20.XA2a.MN0.D a_9848_43396# 7.39e-20
C10201 AVDD a_12368_46916# 0.359f
C10202 XA8.XA1.XA5.MN2.G XA7.XA6.MN2.D 6.33e-19
C10203 a_11000_51140# D<4> 0.0672f
C10204 a_9848_51140# XA4.XA6.MN2.D 0.00176f
C10205 XA0.XA6.MP2.G XA0.XA6.MN2.D 1.59e-19
C10206 XA7.XA9.MN1.G a_18560_50084# 0.00969f
C10207 XA2.XA1.XA5.MN2.G a_2288_50788# 0.00548f
C10208 XA2.XA9.MN1.G a_4808_49732# 0.00119f
C10209 XB1.XA3.MN1.D m3_n1960_4356# 0.0634f
C10210 XA20.XA2a.MN0.D a_8480_40932# 0.0733f
C10211 EN a_12368_42692# 0.159f
C10212 XA2.XA6.MP0.G XA1.XA4.MN0.D 2.8e-19
C10213 D<3> a_12368_48676# 0.00918f
C10214 D<7> a_2288_48324# 0.0164f
C10215 XA20.XA3.MN1.D XA20.XA3.MN0.D 0.547f
C10216 XA8.XA1.XA5.MN2.G XA7.XA4.MN0.G 0.158f
C10217 XA7.XA1.XA5.MN2.G XA8.XA4.MN0.G 3.9e-20
C10218 AVDD a_2288_43748# 0.357f
C10219 XA5.XA6.MN0.D a_13520_49732# 0.00176f
C10220 SARN XA2.XA3.MN0.G 0.0764f
C10221 a_11000_50084# a_12368_50084# 8.89e-19
C10222 SARP a_11000_2446# 0.00767f
C10223 D<8> XDAC2.XC128b<2>.XRES8.B 4.06e-21
C10224 a_n232_42340# a_n232_41988# 0.0109f
C10225 VREF a_9848_47268# 1.19e-19
C10226 XA2.XA6.MP0.G a_4808_46212# 7.76e-20
C10227 XA6.XA6.MP0.G a_16040_46564# 5.5e-19
C10228 a_4808_48324# a_5960_48324# 0.00133f
C10229 XA6.XA1.XA5.MN2.G a_13520_44804# 1.86e-19
C10230 AVDD XA5.XA1.XA1.MN0.S 1.03f
C10231 XA4.XA11.MN1.G XA5.XA11.MN1.G 0.0251f
C10232 AVDD a_22448_53252# 0.388f
C10233 XA4.XA1.XA1.MN0.S a_9848_40228# 0.0215f
C10234 XA4.XA1.XA1.MP1.D a_11000_40932# 0.0465f
C10235 a_23600_41284# a_23600_40932# 0.0109f
C10236 a_7328_46916# a_7328_46564# 0.0109f
C10237 XA7.XA4.MN0.G a_17408_45508# 6.57e-19
C10238 XA2.XA1.XA5.MN2.G a_3440_42340# 4.69e-19
C10239 XA8.XA1.XA5.MN2.G XA8.XA1.XA4.MN0.D 0.00313f
C10240 a_17408_46916# XA7.XA3.MN0.G 0.0674f
C10241 D<8> XA1.XA3.MN0.G 3.29f
C10242 AVDD a_14960_n18# 0.445f
C10243 XA5.XA6.MP0.G XA5.XA1.XA5.MN0.D 7.41e-19
C10244 XA0.XA4.MN0.D EN 0.0648f
C10245 XA1.XA6.MP0.G a_2288_43396# 5.5e-19
C10246 AVDD XA8.XA6.MN2.D 3.58e-19
C10247 CK_SAMPLE a_16040_51140# 8.45e-19
C10248 XA6.XA10.MP0.G a_14888_52548# 0.128f
C10249 a_23600_52900# a_23600_52548# 0.0109f
C10250 XB1.XA1.MP0.D XB1.M1.G 0.129f
C10251 D<2> a_16040_40228# 7.76e-20
C10252 XA20.XA3a.MN0.D a_8480_43044# 0.0905f
C10253 SARN li_14804_31872# 0.00103f
C10254 a_8480_45156# a_9848_45156# 8.89e-19
C10255 XA1.XA1.XA5.MN2.D a_2288_44804# 0.156f
C10256 XA8.XA1.XA5.MN2.D a_19928_45156# 0.153f
C10257 XA5.XA4.MN0.G XA5.XA1.XA4.MN1.D 0.0642f
C10258 D<6> a_5960_39876# 7.76e-20
C10259 XA2.XA9.MN1.G a_4808_50436# 0.01f
C10260 XA20.XA10.MN1.D a_23600_49380# 0.00408f
C10261 AVDD a_n232_47972# 0.00125f
C10262 XA7.XA9.MN1.G a_17408_50788# 0.00281f
C10263 XA4.XA7.MP0.D D<4> 2.65e-19
C10264 XA5.XA11.MP0.D VREF 0.00176f
C10265 XDAC2.XC64b<1>.XRES8.B XDAC2.X16ab.XRES8.B 6.7e-19
C10266 li_14804_27168# li_14804_26556# 0.00271f
C10267 XA0.XA6.MP2.G XDAC1.XC128a<1>.XRES1A.B 0.00406f
C10268 EN XA8.XA1.XA2.MP0.D 0.03f
C10269 XA20.XA3a.MN0.D a_7328_40580# 0.0658f
C10270 XA20.XA2a.MN0.D a_14888_41636# 0.0144f
C10271 SARP a_22448_43044# 5.88e-19
C10272 XA4.XA1.XA5.MP1.D XA4.XA1.XA5.MP0.D 0.0488f
C10273 a_14888_43748# a_16040_43748# 0.00133f
C10274 a_13520_50436# XA5.XA6.MN0.D 0.00176f
C10275 D<7> VREF 1.3f
C10276 XA0.XA6.MP2.G XA3.XA4.MN0.D 0.047f
C10277 AVDD a_13520_44804# 0.00125f
C10278 XA2.XA1.XA5.MN2.G a_2288_49028# 0.00363f
C10279 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES2.B 0.0136f
C10280 XDAC2.XC64a<0>.XRES4.B XDAC2.XC64a<0>.XRES8.B 0.471f
C10281 XA0.XA4.MN0.D li_9184_5676# 0.00506f
C10282 XA1.XA1.XA4.MN1.D a_3440_42340# 0.00176f
C10283 a_16040_42692# a_17408_42692# 8.89e-19
C10284 XA6.XA1.XA5.MN2.G a_12368_45860# 0.00363f
C10285 D<7> a_3440_46212# 0.0141f
C10286 a_23600_49380# a_23600_49028# 0.0109f
C10287 AVDD XA20.XA1.MN0.D 0.478f
C10288 XA2.XA4.MN0.D a_5960_48324# 0.0698f
C10289 AVDD a_19928_53956# 0.00164f
C10290 a_14888_54308# a_16040_54308# 0.00133f
C10291 a_2288_54308# a_2288_53956# 0.0109f
C10292 SARP li_9184_21432# 0.00103f
C10293 a_2288_41284# a_3440_41284# 0.00133f
C10294 XA4.XA6.MP0.G a_9848_44100# 7.76e-20
C10295 XA0.XA6.MP0.G EN 0.0673f
C10296 XA3.XA4.MN0.G a_9848_46564# 2.2e-19
C10297 XA4.XA4.MN0.G a_8480_46564# 2.2e-19
C10298 a_18560_47620# a_18560_47268# 0.0109f
C10299 XA0.XA6.MP2.G a_920_43396# 7.76e-20
C10300 XA4.XA1.XA5.MN2.G a_8480_43044# 2.31e-19
C10301 VREF a_12368_45156# 0.0195f
C10302 XA3.XA4.MN0.D a_8480_45156# 9.24e-20
C10303 AVDD a_9560_2798# 0.00165f
C10304 XA7.XA11.MN1.G XA7.XA9.MN1.G 0.00349f
C10305 XA2.XA10.MP0.D a_5960_52900# 0.0893f
C10306 AVDD a_3440_51492# 0.00166f
C10307 CK_SAMPLE XA8.XA7.MP0.D 0.0217f
C10308 a_12368_39876# a_13520_39876# 0.00133f
C10309 XA2.XA3.MN0.G SARP 0.0395f
C10310 XA7.XA3.MN0.G a_18560_44804# 0.0404f
C10311 D<8> a_920_44452# 0.055f
C10312 XA3.XA4.MN0.G XA3.XA1.XA2.MP0.D 0.206f
C10313 SARN a_9560_2446# 4.94e-19
C10314 XA4.XA1.XA5.MN2.G a_7328_40580# 0.0431f
C10315 XA3.XA1.XA5.MN2.G a_8480_40580# 0.0806f
C10316 XA0.XA6.MP2.G a_n232_40932# 5.24e-19
C10317 XA20.XA3a.MN0.D a_3440_43748# 0.00228f
C10318 a_13520_45860# a_13520_45508# 0.0109f
C10319 XA1.XA9.MN1.G a_2288_51140# 0.0222f
C10320 AVDD a_22448_49380# 0.368f
C10321 a_7328_51844# a_8480_51844# 0.00133f
C10322 XA7.XA7.MP0.D a_18560_51844# 0.159f
C10323 XA1.XA7.MP0.D XA1.XA8.MP0.D 0.124f
C10324 a_18560_52196# XA7.XA8.MP0.D 2.11e-19
C10325 CK_SAMPLE a_19928_49732# 0.0681f
C10326 XA8.XA9.MN1.G a_21080_51492# 6.57e-19
C10327 XA20.XA10.MN1.D XA20.XA3.MN1.D 0.0105f
C10328 a_14888_44100# EN 0.00576f
C10329 XA20.XA2a.MN0.D XA0.XA1.XA4.MN0.D 0.0375f
C10330 D<7> li_9184_27168# 0.00504f
C10331 XA3.XA3.MN0.G a_8480_42340# 0.0029f
C10332 AVDD a_12368_45860# 0.356f
C10333 a_9848_50788# a_11000_50788# 0.00133f
C10334 a_11000_51844# VREF 0.00396f
C10335 XA2.XA1.XA5.MN2.G a_2288_50084# 0.00366f
C10336 EN a_920_41636# 0.00649f
C10337 XA8.XA1.XA2.MP0.D a_21080_42692# 7.68e-20
C10338 XA4.XA1.XA2.MP0.D XA4.XA1.XA4.MP0.D 4.34e-19
C10339 a_7328_43044# XA3.XA1.XA4.MP1.D 0.00176f
C10340 XA2.XA4.MN0.D XA3.XA4.MN0.D 0.935f
C10341 VREF XA5.XA4.MN0.D 0.593f
C10342 XA20.XA3.MN1.D a_23600_49028# 0.0137f
C10343 D<3> a_12368_47620# 0.0147f
C10344 D<7> a_2288_47268# 0.0148f
C10345 XA5.XA1.XA5.MN2.G a_12368_46916# 7.1e-20
C10346 XA6.XA1.XA5.MN2.G a_11000_46916# 7.1e-20
C10347 AVDD a_5960_43044# 0.381f
C10348 a_18560_41988# a_18560_41636# 0.0109f
C10349 XA3.XA1.XA5.MN2.G a_4808_43748# 1.95e-19
C10350 XA8.XA1.XA5.MN2.G XA8.XA1.XA5.MP1.D 5.21e-20
C10351 XA8.XA7.MP0.G XA8.XA1.XA5.MN1.D 6.68e-19
C10352 XA3.XA4.MN0.G a_7328_47620# 0.155f
C10353 VREF a_9848_46212# 7.12e-19
C10354 AVDD a_4808_40580# 0.00125f
C10355 a_12368_47972# a_13520_47972# 0.00133f
C10356 D<1> a_18560_44452# 5.26e-19
C10357 XA2.XA6.MP0.G a_5960_45156# 5.5e-19
C10358 XA5.XA6.MP0.G XA5.XA1.XA5.MN2.D 0.0325f
C10359 a_n232_47972# a_n232_47620# 0.0109f
C10360 D<5> a_8480_44100# 6.49e-19
C10361 XA20.XA10.MN1.D a_22448_53252# 0.0703f
C10362 a_9848_53604# a_9848_53252# 0.0109f
C10363 a_21080_53604# XA8.XA11.MP0.D 0.00176f
C10364 DONE a_22448_52548# 0.00486f
C10365 XA1.XA12.MP0.G a_2288_52900# 1.28e-19
C10366 XA2.XA11.MN1.G a_3440_52900# 0.00295f
C10367 XA6.XA11.MN1.G XA5.XA10.MP0.D 0.0327f
C10368 AVDD XA4.XA9.MN1.G 0.93f
C10369 a_5960_40580# a_5960_40228# 0.0109f
C10370 a_5960_46212# a_7328_46212# 8.89e-19
C10371 a_19928_46564# a_19928_46212# 0.0109f
C10372 D<3> a_12368_41988# 7.77e-20
C10373 D<8> a_920_45508# 0.0698f
C10374 XA7.XA3.MN0.G a_17408_45860# 0.155f
C10375 D<7> a_2288_41636# 7.77e-20
C10376 XA5.XA1.XA5.MN2.G XA5.XA1.XA1.MN0.S 0.0916f
C10377 XA0.XA11.MN1.G a_11000_1038# 0.00151f
C10378 XA7.XA6.MP0.G XA7.XA1.XA4.MP1.D 0.00121f
C10379 XA1.XA4.MN0.D a_2288_43396# 9.15e-20
C10380 XA0.XA4.MN0.G a_n232_44100# 0.0164f
C10381 CK_SAMPLE a_19928_50436# 0.161f
C10382 AVDD XA20.XA3.MN6.D 5.96f
C10383 XA0.XA10.MP0.G XA0.XA8.MP0.D 0.0434f
C10384 XB2.XA3.MN1.D a_14960_1038# 0.0114f
C10385 XB1.XA3.MN1.D a_9560_686# 4.45e-19
C10386 a_11000_1390# a_11000_1038# 0.0109f
C10387 XA5.XA3.MN0.G a_13520_43044# 3.62e-20
C10388 XA3.XA4.MN0.G a_7328_41988# 5.1e-20
C10389 a_3440_45156# EN 4.58e-19
C10390 XA7.XA6.MP0.G a_16040_40228# 5.06e-19
C10391 SARN XDAC2.XC128b<2>.XRES8.B 27.7f
C10392 XA20.XA3a.MN0.D a_n232_42340# 0.00542f
C10393 XA20.XA2a.MN0.D a_8480_43396# 4.8e-20
C10394 a_n232_44452# a_920_44452# 0.00133f
C10395 a_13520_44804# a_13520_44452# 0.0109f
C10396 XA3.XA6.MP0.G a_5960_39876# 1.28e-19
C10397 AVDD a_11000_46916# 0.359f
C10398 XA8.XA1.XA5.MN2.G XA7.XA6.MP2.D 0.00313f
C10399 XA7.XA9.MN1.G a_17408_50084# 0.00281f
C10400 a_7328_52548# VREF 0.00396f
C10401 XA0.XA7.MP0.G a_2288_50788# 7.1e-20
C10402 XA2.XA1.XA5.MN2.G a_920_50788# 7.1e-20
C10403 XB1.XA3.MN1.D m3_n2104_4356# 0.17f
C10404 li_9184_22044# li_9184_21432# 0.00271f
C10405 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES2.B 0.0307f
C10406 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES16.B 0.0381f
C10407 XDAC1.X16ab.XRES1A.B XDAC1.XC128b<2>.XRES1A.B 0.00444f
C10408 XA20.XA2a.MN0.D a_7328_40932# 0.0662f
C10409 XA1.XA1.XA5.MN0.D a_3440_43044# 0.00176f
C10410 XA5.XA1.XA5.MN0.D a_13520_43396# 0.0474f
C10411 a_n232_43396# a_920_43396# 0.00133f
C10412 EN a_11000_42692# 0.159f
C10413 XA20.XA3.MN1.D a_23600_50084# 0.055f
C10414 XA20.XA3.MN6.D XA20.XA3.MN0.D 0.338f
C10415 XA2.XA6.MP0.G VREF 0.568f
C10416 XA8.XA1.XA5.MN2.G XA6.XA4.MN0.G 6.95e-19
C10417 XA7.XA1.XA5.MN2.G XA7.XA4.MN0.G 0.169f
C10418 XA1.XA6.MP0.G XA3.XA4.MN0.D 0.066f
C10419 AVDD a_920_43748# 0.357f
C10420 SARN XA1.XA3.MN0.G 0.137f
C10421 XDAC2.XC1.XRES16.B li_14804_6288# 0.00117f
C10422 XDAC1.XC1.XRES16.B XDAC1.XC1.XRES1A.B 0.454f
C10423 SARP a_9560_2446# 0.00101f
C10424 XA4.XA1.XA4.MP0.D a_11000_41988# 0.00176f
C10425 a_11000_42340# a_12368_42340# 8.89e-19
C10426 XA6.XA6.MP0.G a_14888_46564# 5e-19
C10427 a_17408_48676# a_17408_48324# 0.0109f
C10428 D<4> XA4.XA1.XA5.MN2.D 0.0347f
C10429 XA6.XA1.XA5.MN2.G a_12368_44804# 0.00486f
C10430 XA5.XA1.XA5.MN2.G a_13520_44804# 1.95e-19
C10431 D<1> a_18560_45508# 0.0031f
C10432 XA20.XA10.MN1.D XA20.XA1.MN0.D 0.112f
C10433 AVDD XA4.XA1.XA1.MP2.D 0.127f
C10434 XA2.XA4.MN0.D a_5960_47268# 0.0576f
C10435 VREF a_8480_47268# 1.19e-19
C10436 XA3.XA11.MN1.G XA4.XA12.MP0.G 0.00122f
C10437 XA4.XA11.MN1.G XA3.XA12.MP0.G 0.391f
C10438 a_8480_53956# a_8480_53604# 0.0109f
C10439 AVDD a_21080_53252# 0.364f
C10440 a_21080_53956# XA8.XA12.MP0.G 0.0658f
C10441 XA4.XA1.XA1.MN0.D a_11000_40932# 8.29e-20
C10442 SARP XDAC1.XC64a<0>.XRES8.B 27.7f
C10443 XA0.XA4.MN0.G XA0.XA1.XA5.MN2.D 0.135f
C10444 XA2.XA1.XA5.MN2.G a_2288_42340# 0.00442f
C10445 XA0.XA7.MP0.G a_3440_42340# 0.00568f
C10446 XA8.XA1.XA5.MN2.G XA7.XA1.XA4.MN0.D 7.72e-19
C10447 AVDD a_13808_n18# 0.00236f
C10448 D<2> XA6.XA1.XA4.MP1.D 7.42e-19
C10449 XA5.XA6.MP0.G XA5.XA1.XA5.MP0.D 0.00121f
C10450 CK_SAMPLE a_14888_51140# 0.0686f
C10451 a_3440_52548# a_4808_52548# 8.89e-19
C10452 XA20.XA9.MP0.D SARN 0.652f
C10453 AVDD D<0> 2.26f
C10454 D<2> a_14888_40228# 6.49e-19
C10455 XA20.XA3a.MN0.D a_7328_43044# 0.00877f
C10456 XA5.XA4.MN0.G XA5.XA1.XA4.MP1.D 0.0488f
C10457 XA4.XA3.MN0.G a_9848_43748# 2.78e-19
C10458 D<6> a_4808_39876# 0.00197f
C10459 XA2.XA4.MN0.D a_5960_41636# 9.14e-20
C10460 XA20.XA10.MN1.D a_22448_49380# 1.69e-19
C10461 AVDD XA8.XA4.MN0.G 2.39f
C10462 CK_SAMPLE a_19928_48676# 1.95e-19
C10463 a_5960_51492# XA3.XA1.XA5.MN2.G 0.0699f
C10464 a_17408_52196# D<1> 7.56e-20
C10465 a_16040_51492# a_17408_51492# 8.89e-19
C10466 XA4.XA11.MP0.D VREF 0.00185f
C10467 EN XA7.XA1.XA5.MN0.D 0.0063f
C10468 XA20.XA3a.MN0.D a_5960_40580# 0.0674f
C10469 XA20.XA2a.MN0.D a_13520_41636# 0.0145f
C10470 XA0.XA6.MP2.D VREF 5.13e-19
C10471 XA0.XA6.MP2.G XA2.XA4.MN0.D 0.0481f
C10472 D<7> XA0.XA4.MN0.D 2.87f
C10473 XA1.XA6.MP0.G XA1.XA6.MP0.D 0.0392f
C10474 AVDD a_12368_44804# 0.356f
C10475 XA20.XA9.MP0.D a_23600_46916# 0.00334f
C10476 XA0.XA7.MP0.G a_2288_49028# 7.1e-20
C10477 XA2.XA1.XA5.MN2.G a_920_49028# 7.1e-20
C10478 XA6.XA1.XA4.MN1.D XA6.XA1.XA4.MN0.D 0.0488f
C10479 a_3440_42692# XA1.XA1.XA4.MN0.D 0.00176f
C10480 D<8> XDAC2.XC0.XRES8.B 0.00688f
C10481 XA6.XA1.XA5.MN2.G a_11000_45860# 7.1e-20
C10482 XA5.XA1.XA5.MN2.G a_12368_45860# 7.1e-20
C10483 D<7> a_2288_46212# 0.0202f
C10484 D<6> XA20.XA2a.MN0.D 0.0752f
C10485 a_9848_49028# a_11000_49028# 0.00133f
C10486 AVDD XA8.XA1.XA4.MP0.D 0.147f
C10487 VREF a_7328_48324# 0.0536f
C10488 XA2.XA4.MN0.D a_4808_48324# 0.0981f
C10489 D<3> a_13520_46564# 0.0551f
C10490 AVDD a_18560_53956# 0.00166f
C10491 XA0.XA1.XA1.MP2.D XA0.XA1.XA1.MP1.D 0.0488f
C10492 XA3.XA4.MN0.G a_8480_46564# 0.0155f
C10493 a_4808_47268# a_5960_47268# 0.00133f
C10494 XA0.XA6.MP2.G a_n232_43396# 6.49e-19
C10495 XA3.XA1.XA5.MN2.G a_8480_43044# 0.0732f
C10496 XA4.XA1.XA5.MN2.G a_7328_43044# 0.00551f
C10497 VREF a_11000_45156# 0.0195f
C10498 XA3.XA4.MN0.D a_7328_45156# 9.15e-20
C10499 AVDD a_8408_2798# 0.464f
C10500 XA6.XA12.MP0.G XA6.XA9.MN1.G 4.5e-19
C10501 a_16040_53252# a_16040_52900# 0.0109f
C10502 XA2.XA10.MP0.D a_4808_52900# 0.128f
C10503 AVDD a_2288_51492# 0.387f
C10504 CK_SAMPLE XA7.XA7.MP0.D 0.00428f
C10505 XA1.XA3.MN0.G SARP 0.0622f
C10506 XA7.XA3.MN0.G a_17408_44804# 0.00498f
C10507 D<8> a_n232_44452# 0.096f
C10508 XA3.XA1.XA5.MN2.G a_7328_40580# 0.00417f
C10509 XA20.XA3a.MN0.D a_2288_43748# 0.00106f
C10510 a_920_45860# XA0.XA1.XA5.MN2.D 3.12e-20
C10511 a_n232_45508# a_920_45508# 0.00133f
C10512 AVDD a_21080_49380# 0.356f
C10513 XA7.XA7.MP0.D a_17408_51844# 0.133f
C10514 a_17408_54308# VREF 0.00579f
C10515 CK_SAMPLE a_18560_49732# 0.0709f
C10516 XA8.XA9.MN1.G a_19928_51492# 0.0118f
C10517 XA20.XA10.MN1.D XA20.XA3.MN6.D 0.196f
C10518 XA4.XA9.MN1.G XA5.XA1.XA5.MN2.G 0.0494f
C10519 XDAC1.XC0.XRES8.B li_9184_31872# 9.91e-20
C10520 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES16.B 0.0381f
C10521 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES2.B 0.0307f
C10522 li_14804_32484# li_14804_31872# 0.00271f
C10523 a_5960_44100# XA2.XA1.XA5.MP1.D 0.00176f
C10524 a_13520_44100# EN 0.00576f
C10525 a_18560_44100# a_19928_44100# 8.89e-19
C10526 XA20.XA3a.MN0.D XA5.XA1.XA1.MN0.S 0.0673f
C10527 XA5.XA1.XA5.MN2.D a_13520_43396# 1.28e-19
C10528 XA20.XA2a.MN0.D a_23600_42692# 0.00306f
C10529 XA0.XA6.MP2.G XDAC1.XC64b<1>.XRES1A.B 4.06e-21
C10530 SARN li_14804_11604# 0.00103f
C10531 AVDD a_11000_45860# 0.356f
C10532 XA8.XA6.MP2.D a_21080_50788# 0.049f
C10533 XA2.XA1.XA5.MN2.G a_920_50084# 7.1e-20
C10534 XA0.XA7.MP0.G a_2288_50084# 7.1e-20
C10535 D<7> XA0.XA6.MP0.G 0.0688f
C10536 XA4.XA6.MP2.D a_11000_50436# 0.00176f
C10537 XA8.XA7.MP0.G XA8.XA6.MP0.G 0.042f
C10538 XDAC2.XC128a<1>.XRES16.B XDAC2.XC128a<1>.XRES1A.B 0.454f
C10539 EN a_n232_41636# 0.00426f
C10540 XA20.XA2a.MN0.D a_19928_39876# 1.09e-19
C10541 XA4.XA1.XA2.MP0.D XA4.XA1.XA4.MN0.D 0.056f
C10542 XA0.XA1.XA2.MP0.D a_920_42340# 2.54e-19
C10543 XA8.XA1.XA2.MP0.D a_19928_42692# 0.0962f
C10544 a_18560_43044# a_19928_43044# 8.89e-19
C10545 XA0.XA6.MP0.G XDAC2.XC1.XRES1A.B 0.00405f
C10546 XA20.XA3.MN6.D a_23600_49028# 5.18e-19
C10547 a_21080_49732# XA8.XA4.MN0.D 0.0658f
C10548 VREF XA4.XA4.MN0.D 0.593f
C10549 XA20.XA3.MN1.D a_22448_49028# 0.00253f
C10550 XA1.XA4.MN0.D XA3.XA4.MN0.D 0.0357f
C10551 XA20.XA9.MP0.D SARP 0.405f
C10552 XA5.XA1.XA5.MN2.G a_11000_46916# 0.00455f
C10553 AVDD a_4808_43044# 0.00125f
C10554 a_9848_49732# a_9848_49380# 0.0109f
C10555 a_5960_41988# XA2.XA1.XA1.MN0.S 3.8e-19
C10556 a_4808_41636# a_5960_41636# 0.00133f
C10557 SARP li_9184_31872# 0.00103f
C10558 VREF a_8480_46212# 7.12e-19
C10559 XA2.XA4.MN0.D a_5960_46212# 9.14e-20
C10560 XA2.XA1.XA5.MN2.G a_4808_43748# 0.0732f
C10561 XA8.XA1.XA5.MN2.G XA8.XA1.XA5.MN1.D 0.0102f
C10562 AVDD a_3440_40580# 0.00125f
C10563 D<1> a_17408_44452# 1.48e-19
C10564 XA2.XA6.MP0.G a_4808_45156# 7.76e-20
C10565 D<5> a_7328_44100# 7.77e-20
C10566 DONE a_21080_52548# 0.00228f
C10567 AVDD XA3.XA9.MN0.D 4.25e-19
C10568 XA2.XA11.MN1.G a_2288_52900# 1.34e-19
C10569 a_17408_40580# a_18560_40580# 0.00133f
C10570 XA20.XA3a.MN0.D a_13520_44804# 1.57e-20
C10571 XA3.XA6.MP0.G a_8480_42692# 7.76e-20
C10572 D<8> a_n232_45508# 0.107f
C10573 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MP2.D 0.0736f
C10574 XA6.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S 3.84e-21
C10575 XA0.XA11.MN1.G a_9560_1038# 0.00173f
C10576 VREF a_2288_43396# 3.39e-19
C10577 XA6.XA4.MN0.G a_16040_44452# 5.54e-19
C10578 CK_SAMPLE a_18560_50436# 0.161f
C10579 XA20.XA10.MN1.D D<0> 0.00217f
C10580 AVDD XA20.XA3a.MN0.G 5.77f
C10581 a_14888_52548# XA6.XA7.MP0.D 5.16e-20
C10582 a_23600_52548# a_23600_52196# 0.0109f
C10583 XA6.XA10.MP0.G a_16040_51844# 0.00224f
C10584 XB1.XA3.MN0.S a_9560_686# 0.0328f
C10585 XB1.XA3.MN1.D a_8408_686# 0.00656f
C10586 XB2.XA3.MN0.S a_14960_1038# 0.00224f
C10587 XB2.XA3.MN1.D a_13808_1038# 0.00252f
C10588 a_13808_1390# a_14960_1390# 0.00133f
C10589 XA7.XA6.MP0.G a_14888_40228# 7.45e-19
C10590 a_2288_45156# EN 1.83e-19
C10591 XA3.XA1.XA5.MN2.D XA3.XA1.XA5.MN1.D 0.0488f
C10592 XA0.XA7.MP0.G a_920_50788# 0.00548f
C10593 AVDD a_9848_46916# 0.00131f
C10594 XA8.XA1.XA5.MN2.G D<1> 0.704f
C10595 a_5960_52548# VREF 0.00396f
C10596 XB1.XA3.MN1.D m3_7544_4532# 0.0137f
C10597 XA20.XA2a.MN0.D a_5960_40932# 0.0678f
C10598 XA5.XA1.XA5.MN0.D a_12368_43396# 2.16e-19
C10599 XA5.XA1.XA5.MP0.D a_13520_43396# 2.16e-19
C10600 XA20.XA3.MN6.D a_23600_50084# 0.00276f
C10601 XA20.XA3a.MN0.G XA20.XA3.MN0.D 0.357f
C10602 XA2.XA1.XA5.MN2.G a_2288_47972# 0.00363f
C10603 XA5.XA6.MP0.D a_12368_49732# 0.00176f
C10604 XA5.XA6.MP0.G a_13520_49732# 0.00239f
C10605 XA2.XA6.MP0.G XA0.XA4.MN0.D 1.9e-19
C10606 XA7.XA1.XA5.MN2.G XA6.XA4.MN0.G 0.158f
C10607 XA20.XA9.MP0.D a_23600_45860# 0.00334f
C10608 XA1.XA6.MP0.G XA2.XA4.MN0.D 0.0732f
C10609 AVDD a_n232_43748# 0.00125f
C10610 SARN D<8> 0.327f
C10611 a_9848_50084# a_11000_50084# 0.00133f
C10612 D<8> li_14804_22044# 3.5e-20
C10613 XA20.XA1.MN0.D a_23600_42340# 0.0529f
C10614 XA3.XA6.MP0.G XA20.XA2a.MN0.D 0.0699f
C10615 a_3440_48324# a_4808_48324# 8.89e-19
C10616 D<7> a_3440_45156# 7.77e-19
C10617 XA5.XA1.XA5.MN2.G a_12368_44804# 7.1e-20
C10618 XA6.XA1.XA5.MN2.G a_11000_44804# 7.1e-20
C10619 D<1> a_17408_45508# 0.00436f
C10620 AVDD XA4.XA1.XA1.MN0.S 1.04f
C10621 VREF a_7328_47268# 0.0191f
C10622 XA2.XA4.MN0.D a_4808_47268# 0.0963f
C10623 XA2.XA12.MP0.G XA3.XA12.MP0.G 0.00217f
C10624 AVDD a_19928_53252# 0.00154f
C10625 a_19928_53956# XA8.XA12.MP0.G 0.0704f
C10626 XA4.XA1.XA1.MN0.D a_9848_40932# 0.0535f
C10627 a_22448_41284# a_22448_40932# 0.0109f
C10628 a_5960_46916# a_5960_46564# 0.0109f
C10629 XA0.XA7.MP0.G a_2288_42340# 1.97e-19
C10630 XA7.XA1.XA5.MN2.G XA7.XA1.XA4.MN0.D 0.00313f
C10631 XA8.XA1.XA5.MN2.G XA7.XA1.XA4.MP0.D 0.00361f
C10632 a_16040_46916# XA6.XA3.MN0.G 0.0658f
C10633 AVDD a_12368_n18# 7e-19
C10634 D<2> XA6.XA1.XA4.MN1.D 0.00188f
C10635 XA5.XA6.MP0.G XA5.XA1.XA2.MP0.D 0.0125f
C10636 VREF a_21080_44100# 0.0251f
C10637 XA6.XA4.MN0.G a_16040_45508# 6.57e-19
C10638 AVDD XA7.XA6.MN2.D 3.77e-19
C10639 CK_SAMPLE a_13520_51140# 0.067f
C10640 XA5.XA10.MP0.G a_13520_52548# 0.13f
C10641 a_22448_52900# a_22448_52548# 0.0109f
C10642 a_9848_52900# XA4.XA9.MN1.G 0.00113f
C10643 SAR_IP a_11000_2446# 0.0495f
C10644 a_14960_2798# a_14960_2446# 0.0109f
C10645 a_14960_3150# XB2.XA4.MP0.D 0.00252f
C10646 XA20.XA3a.MN0.D a_5960_43044# 0.00835f
C10647 SARN XDAC2.XC0.XRES8.B 27.7f
C10648 a_7328_45156# a_8480_45156# 0.00133f
C10649 XA0.XA1.XA5.MN2.D a_920_44804# 0.156f
C10650 XA7.XA1.XA5.MN2.D a_18560_45156# 0.153f
C10651 XA3.XA3.MN0.G a_9848_43748# 7.98e-19
C10652 XA4.XA6.MP0.G XA4.XA1.XA1.MN0.D 0.00159f
C10653 XA2.XA4.MN0.D a_4808_41636# 9.25e-20
C10654 AVDD XA7.XA4.MN0.G 2.36f
C10655 CK_SAMPLE a_18560_48676# 4.46e-19
C10656 a_2288_51844# D<7> 1.25e-19
C10657 a_4808_51492# XA3.XA1.XA5.MN2.G 0.0674f
C10658 XA3.XA11.MP0.D VREF 0.00176f
C10659 XDAC1.XC64b<1>.XRES8.B XDAC1.X16ab.XRES8.B 6.7e-19
C10660 li_9184_27168# li_9184_26556# 0.00271f
C10661 XA0.XA6.MP2.G li_9184_16728# 0.00508f
C10662 EN XA7.XA1.XA5.MP0.D 0.0446f
C10663 XA2.XA6.MP0.G XDAC2.XC64b<1>.XRES16.B 2.19e-20
C10664 XA20.XA3a.MN0.D a_4808_40580# 0.0658f
C10665 XA20.XA2a.MN0.D a_12368_41636# 0.00184f
C10666 XA4.XA1.XA5.MP1.D XA4.XA1.XA2.MP0.D 6.52e-20
C10667 XA4.XA1.XA5.MN1.D XA4.XA1.XA5.MN0.D 0.0488f
C10668 a_13520_43748# a_14888_43748# 8.89e-19
C10669 a_920_43748# XA0.XA1.XA5.MP0.D 0.00176f
C10670 XA0.XA6.MP2.G XA1.XA4.MN0.D 0.0101f
C10671 a_22448_50788# XA20.XA3.MN6.D 1.06e-19
C10672 XA0.XA6.MP0.G XA2.XA6.MP0.G 0.0722f
C10673 XA8.XA1.XA5.MN2.G a_17408_49380# 0.00363f
C10674 a_13520_50436# XA5.XA6.MP0.G 3.02e-20
C10675 a_12368_50436# XA5.XA6.MP0.D 0.00176f
C10676 AVDD a_11000_44804# 0.356f
C10677 XA0.XA7.MP0.G a_920_49028# 0.00363f
C10678 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES2.B 0.0136f
C10679 XDAC1.XC64a<0>.XRES4.B XDAC1.XC64a<0>.XRES8.B 0.471f
C10680 XA0.XA4.MN0.D XDAC1.XC1.XRES1A.B 0.00405f
C10681 XA6.XA1.XA2.MP0.D a_16040_41636# 0.00224f
C10682 XA1.XA1.XA4.MP1.D a_2288_42340# 0.00176f
C10683 a_14888_42692# a_16040_42692# 0.00133f
C10684 D<8> XDAC1.XC0.XRES8.B 7.76e-19
C10685 a_22448_49380# a_22448_49028# 0.0109f
C10686 XA5.XA1.XA5.MN2.G a_11000_45860# 0.00363f
C10687 AVDD XA8.XA1.XA4.MN0.D 0.00913f
C10688 VREF a_5960_48324# 0.0536f
C10689 XA8.XA4.MN0.D a_21080_48676# 0.154f
C10690 XA20.XA3.MN6.D XA20.XA3a.MN0.D 0.449f
C10691 D<3> a_12368_46564# 0.0695f
C10692 AVDD a_17408_53956# 0.464f
C10693 a_13520_54308# a_14888_54308# 8.89e-19
C10694 a_920_54308# a_920_53956# 0.0109f
C10695 SARP XDAC1.XC128b<2>.XRES8.B 27.7f
C10696 XA0.XA1.XA1.MN0.S XA0.XA1.XA1.MP1.D 0.0615f
C10697 XA5.XA1.XA1.MP2.D a_12368_41284# 0.0465f
C10698 a_920_41284# a_2288_41284# 8.89e-19
C10699 XA5.XA1.XA1.MN0.S a_13520_41284# 0.0674f
C10700 XA3.XA4.MN0.G a_7328_46564# 3.46e-19
C10701 a_17408_47620# a_17408_47268# 0.0109f
C10702 D<4> XA4.XA1.XA5.MP0.D 7.42e-19
C10703 VREF a_9848_45156# 7.39e-19
C10704 AVDD a_14960_3150# 0.485f
C10705 DONE a_23600_51844# 1.97e-19
C10706 XA7.XA11.MN1.G XA6.XA9.MN1.G 0.00116f
C10707 XA2.XA11.MN1.G a_3440_52196# 1.84e-19
C10708 XA7.XA10.MP0.D XA8.XA10.MP0.D 0.00217f
C10709 AVDD a_920_51492# 0.387f
C10710 CK_SAMPLE XA6.XA7.MP0.D 0.00417f
C10711 a_11000_39876# a_12368_39876# 8.89e-19
C10712 D<8> SARP 0.2f
C10713 XA2.XA4.MN0.G XA2.XA1.XA5.MP0.D 0.00138f
C10714 D<1> a_18560_41284# 6.49e-19
C10715 XA3.XA1.XA5.MN2.G a_5960_40580# 0.0506f
C10716 D<5> XA3.XA1.XA1.MN0.D 0.0166f
C10717 XA20.XA3a.MN0.D a_920_43748# 0.00106f
C10718 a_12368_45860# a_12368_45508# 0.0109f
C10719 SARN XB2.XA1.MP0.D 0.00571f
C10720 AVDD a_19928_49380# 0.00159f
C10721 a_5960_51844# a_7328_51844# 8.89e-19
C10722 XA0.XA7.MP0.D XA0.XA8.MP0.D 0.124f
C10723 a_16040_54308# VREF 0.00579f
C10724 CK_SAMPLE a_17408_49732# 0.00347f
C10725 XA8.XA9.MN1.G a_18560_51492# 2.84e-19
C10726 XA20.XA10.MN1.D XA20.XA3a.MN0.G 0.15f
C10727 XA4.XA9.MN1.G XA4.XA1.XA5.MN2.G 4.35e-19
C10728 D<7> XDAC1.XC64b<1>.XRES16.B 0.0282f
C10729 a_12368_44100# EN 0.0767f
C10730 XA5.XA1.XA5.MN2.D a_12368_43396# 4.58e-19
C10731 XA20.XA2a.MN0.D a_22448_42692# 0.00611f
C10732 XA0.XA6.MP2.G XA0.XA6.MP0.D 0.0323f
C10733 AVDD a_9848_45860# 0.00125f
C10734 a_8480_50788# a_9848_50788# 8.89e-19
C10735 XA0.XA7.MP0.G a_920_50084# 0.00366f
C10736 XA20.XA2a.MN0.D a_18560_39876# 1.09e-19
C10737 XA0.XA1.XA2.MP0.D a_n232_42340# 0.095f
C10738 a_5960_43044# XA2.XA1.XA4.MP1.D 0.00176f
C10739 a_19928_49732# XA8.XA4.MN0.D 0.0675f
C10740 XA1.XA4.MN0.D XA2.XA4.MN0.D 1.55f
C10741 VREF XA3.XA4.MN0.D 0.615f
C10742 XA20.XA3.MN6.D a_22448_49028# 0.0125f
C10743 XA5.XA6.MP0.G a_13520_48676# 0.0651f
C10744 D<0> XA20.XA3a.MN0.D 2.09e-20
C10745 XA1.XA6.MP0.G a_3440_48324# 0.00295f
C10746 XA20.XA9.MP0.D a_23600_44804# 0.00558f
C10747 AVDD a_3440_43044# 0.00125f
C10748 a_17408_42340# XA7.XA1.XA1.MN0.S 1.34e-19
C10749 a_17408_41988# a_17408_41636# 0.0109f
C10750 XA2.XA4.MN0.D a_4808_46212# 6.37e-19
C10751 VREF a_7328_46212# 0.0671f
C10752 XA2.XA1.XA5.MN2.G a_3440_43748# 2.66e-19
C10753 XA0.XA7.MP0.G a_4808_43748# 7.1e-20
C10754 XA8.XA1.XA5.MN2.G XA7.XA1.XA5.MN1.D 6.68e-19
C10755 XA2.XA4.MN0.G a_5960_47620# 0.155f
C10756 AVDD a_2288_40580# 0.381f
C10757 a_11000_47972# a_12368_47972# 8.89e-19
C10758 XA8.XA4.MN0.G XA20.XA3a.MN0.D 0.0979f
C10759 XA8.XA12.MP0.G a_21080_53252# 0.00276f
C10760 XA0.XA12.MP0.D a_3440_52900# 0.00208f
C10761 XA5.XA11.MN1.G XA5.XA10.MP0.D 0.0909f
C10762 XA4.XA12.MP0.G XA4.XA10.MP0.D 0.0632f
C10763 a_8480_53604# a_8480_53252# 0.0109f
C10764 DONE a_19928_52548# 1.98e-19
C10765 AVDD XA3.XA9.MN1.G 0.93f
C10766 a_4808_40580# a_4808_40228# 0.0109f
C10767 a_18560_46564# a_18560_46212# 0.0109f
C10768 a_4808_46212# a_5960_46212# 0.00133f
C10769 XA3.XA6.MP0.G a_7328_42692# 5.5e-19
C10770 XA6.XA3.MN0.G a_16040_45860# 0.155f
C10771 XA5.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S 0.327f
C10772 VREF a_920_43396# 3.39e-19
C10773 XA6.XA4.MN0.G a_14888_44452# 0.00907f
C10774 CK_SAMPLE a_17408_50436# 0.00312f
C10775 AVDD XA8.XA6.MP0.D 0.157f
C10776 XA6.XA10.MP0.G a_14888_51844# 5.59e-19
C10777 XA4.XA9.MN1.G a_11000_52196# 0.0681f
C10778 XA4.XA9.MN0.D a_9848_52196# 0.0492f
C10779 XB1.XA0.MP0.D a_9560_334# 0.00401f
C10780 XB1.XA3.MN0.S a_8408_686# 0.0215f
C10781 XB2.XA3.MN0.S a_13808_1038# 0.0288f
C10782 a_9560_1390# a_9560_1038# 0.0109f
C10783 SARN li_14804_22044# 0.00103f
C10784 XA0.XA4.MN0.D a_920_40932# 9.14e-20
C10785 XA7.XA6.MP0.G a_13520_40228# 5.06e-19
C10786 a_920_45156# EN 1.83e-19
C10787 XA2.XA6.MP0.G a_7328_39876# 1.28e-19
C10788 XA20.XA3a.MN0.D XA8.XA1.XA4.MP0.D 1.13e-19
C10789 XA3.XA1.XA5.MN2.D XA3.XA1.XA5.MP1.D 0.0488f
C10790 a_12368_44804# a_12368_44452# 0.0109f
C10791 XA2.XA4.MN0.G a_5960_41988# 5.1e-20
C10792 XA0.XA7.MP0.G a_n232_50788# 1.87e-19
C10793 AVDD a_8480_46916# 0.00131f
C10794 a_8480_51140# XA3.XA6.MN2.D 0.00176f
C10795 XA1.XA9.MN1.G a_3440_49732# 0.00119f
C10796 XA7.XA1.XA5.MN2.G D<1> 0.0801f
C10797 XB1.XA3.MN1.D m3_7472_4532# 0.0137f
C10798 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES2.B 0.0136f
C10799 XDAC2.XC128b<2>.XRES4.B XDAC2.XC128b<2>.XRES8.B 0.471f
C10800 XA20.XA2a.MN0.D a_4808_40932# 0.0717f
C10801 XA1.XA1.XA2.MP0.D a_3440_43044# 0.0292f
C10802 XA1.XA1.XA5.MP0.D a_2288_43044# 0.00176f
C10803 XA5.XA1.XA5.MP0.D a_12368_43396# 0.049f
C10804 XA5.XA1.XA2.MP0.D a_13520_43396# 0.0961f
C10805 XA20.XA3.MN6.D a_22448_50084# 0.0631f
C10806 XA20.XA3a.MN0.G a_23600_50084# 0.0674f
C10807 XA2.XA1.XA5.MN2.G a_920_47972# 7.1e-20
C10808 XA0.XA7.MP0.G a_2288_47972# 7.1e-20
C10809 XA5.XA6.MP0.G a_12368_49732# 0.099f
C10810 XA6.XA1.XA5.MN2.G XA6.XA4.MN0.G 0.168f
C10811 XA1.XA6.MP0.G XA1.XA4.MN0.D 4.65f
C10812 XA1.XA6.MP0.D VREF 0.0115f
C10813 AVDD XA8.XA1.XA5.MP1.D 0.0846f
C10814 SARN a_23600_46916# 0.0017f
C10815 XDAC1.XC1.XRES16.B li_9184_6288# 0.00117f
C10816 li_14804_6900# li_14804_6288# 0.00271f
C10817 XDAC2.XC1.XRES2.B XDAC2.XC1.XRES1A.B 0.0136f
C10818 SARP XB2.XA1.MP0.D 0.00453f
C10819 XA20.XA1.MN0.D a_22448_42340# 2.16e-19
C10820 XA5.XA1.XA2.MP0.D a_12368_40932# 4.25e-20
C10821 XA4.XA1.XA4.MN0.D a_9848_41988# 0.00176f
C10822 a_9848_42340# a_11000_42340# 0.00133f
C10823 a_16040_48676# a_16040_48324# 0.0109f
C10824 a_4808_48676# XA2.XA4.MN0.G 1.34e-19
C10825 D<7> a_2288_45156# 6.68e-19
C10826 XA5.XA1.XA5.MN2.G a_11000_44804# 0.00486f
C10827 AVDD XA3.XA1.XA1.MP2.D 0.127f
C10828 VREF a_5960_47268# 0.0191f
C10829 XA8.XA4.MN0.D a_21080_47620# 0.00498f
C10830 XA1.XA4.MN0.D a_4808_47268# 4.76e-20
C10831 XA2.XA4.MN0.D a_3440_47268# 4.76e-20
C10832 a_7328_53956# a_7328_53604# 0.0109f
C10833 XA2.XA12.MP0.G XA4.XA11.MN1.G 1.54e-19
C10834 XA3.XA11.MN1.G XA3.XA12.MP0.G 0.278f
C10835 AVDD a_18560_53252# 0.00144f
C10836 SARP li_9184_11604# 0.00103f
C10837 XA3.XA1.XA1.MN0.S a_8480_40228# 0.0215f
C10838 XA8.XA1.XA1.MN0.S a_21080_40580# 0.0318f
C10839 XA0.XA7.MP0.G a_920_42340# 0.00442f
C10840 XA7.XA1.XA5.MN2.G XA7.XA1.XA4.MP0.D 6.33e-19
C10841 D<6> a_5960_42692# 7.76e-20
C10842 a_14888_46916# XA6.XA3.MN0.G 0.0682f
C10843 AVDD a_11000_n18# 7e-19
C10844 XA6.XA4.MN0.G a_14888_45508# 0.0104f
C10845 a_2288_52548# a_3440_52548# 0.00133f
C10846 XA5.XA10.MP0.G a_12368_52548# 0.0684f
C10847 AVDD XA7.XA6.MP2.D 0.172f
C10848 CK_SAMPLE a_12368_51140# 8.45e-19
C10849 SAR_IN XB2.XA1.MP0.D 0.0168f
C10850 SAR_IP a_9560_2446# 1.82e-19
C10851 XA0.XA6.MP0.G a_920_40932# 4.24e-19
C10852 XA7.XA1.XA5.MN2.D a_17408_45156# 0.155f
C10853 XA0.XA1.XA5.MN2.D a_n232_44804# 0.153f
C10854 XA20.XA3a.MN0.D a_4808_43044# 0.0864f
C10855 XA4.XA4.MN0.G XA4.XA1.XA4.MP1.D 0.0488f
C10856 XA3.XA3.MN0.G a_8480_43748# 0.00371f
C10857 XA20.XA2a.MN0.D EN 0.897f
C10858 AVDD XA6.XA4.MN0.G 2.36f
C10859 CK_SAMPLE a_17408_48676# 6.2e-20
C10860 XA6.XA9.MN1.G a_16040_50788# 0.00281f
C10861 a_14888_51492# a_16040_51492# 0.00133f
C10862 XA2.XA11.MP0.D VREF 0.00185f
C10863 XA1.XA9.MN1.G a_3440_50436# 0.01f
C10864 D<8> a_n232_41284# 0.00335f
C10865 EN XA7.XA1.XA2.MP0.D 0.03f
C10866 XA20.XA3a.MN0.D a_3440_40580# 0.0674f
C10867 XA20.XA2a.MN0.D a_11000_41636# 0.00184f
C10868 XA4.XA1.XA5.MN1.D XA4.XA1.XA2.MP0.D 0.0102f
C10869 D<4> a_11000_49732# 0.0109f
C10870 XA0.XA6.MP2.G VREF 1.3f
C10871 a_22448_50788# XA20.XA3a.MN0.G 6.76e-20
C10872 XA7.XA1.XA5.MN2.G a_17408_49380# 7.1e-20
C10873 XA8.XA1.XA5.MN2.G a_16040_49380# 7.1e-20
C10874 a_12368_50436# XA5.XA6.MP0.G 0.0678f
C10875 AVDD a_9848_44804# 0.00125f
C10876 XA5.XA1.XA4.MN1.D XA5.XA1.XA4.MN0.D 0.0488f
C10877 XA2.XA1.XA2.MP0.D XA2.XA1.XA1.MN0.S 2.11e-19
C10878 XA6.XA1.XA2.MP0.D a_14888_41636# 0.00316f
C10879 a_2288_42692# XA1.XA1.XA4.MP0.D 0.00176f
C10880 D<8> li_14804_32484# 0.00508f
C10881 a_8480_49028# a_9848_49028# 8.89e-19
C10882 XA1.XA6.MP0.G a_3440_47268# 1.38e-19
C10883 AVDD XA7.XA1.XA4.MN0.D 0.00889f
C10884 XA1.XA4.MN0.D a_3440_48324# 0.0997f
C10885 XA8.XA4.MN0.D a_19928_48676# 0.158f
C10886 XA20.XA3a.MN0.G XA20.XA3a.MN0.D 0.515f
C10887 XA20.XA3.MN6.D a_23600_47972# 6.5e-19
C10888 SARN SARP 6.26f
C10889 XA5.XA6.MP0.G a_13520_47620# 4.4e-19
C10890 AVDD a_16040_53956# 0.461f
C10891 XA0.XA1.XA1.MN0.S XA0.XA1.XA1.MN0.D 0.0743f
C10892 XA5.XA1.XA1.MN0.S a_12368_41284# 0.0948f
C10893 a_3440_47268# a_4808_47268# 8.89e-19
C10894 XA3.XA1.XA5.MN2.G a_5960_43044# 0.00551f
C10895 D<4> XA4.XA1.XA5.MN0.D 0.00188f
C10896 XA2.XA4.MN0.D a_5960_45156# 9.14e-20
C10897 VREF a_8480_45156# 7.39e-19
C10898 AVDD a_13808_3150# 0.00166f
C10899 DONE a_22448_51844# 0.00486f
C10900 a_14888_53252# a_14888_52900# 0.0109f
C10901 XA1.XA10.MP0.D a_3440_52900# 0.13f
C10902 AVDD a_n232_51492# 0.00166f
C10903 CK_SAMPLE XA5.XA7.MP0.D 0.00428f
C10904 a_23600_40228# a_23600_39876# 0.0109f
C10905 XA2.XA1.XA5.MN2.G a_5960_40580# 5.68e-19
C10906 D<1> a_17408_41284# 7.77e-20
C10907 XA3.XA1.XA5.MN2.G a_4808_40580# 9.75e-19
C10908 XA8.XA7.MP0.G a_22448_40932# 9.75e-19
C10909 XA5.XA6.MP0.G a_13520_41988# 7.76e-20
C10910 XA20.XA3a.MN0.D a_n232_43748# 0.00218f
C10911 SARN SAR_IN 1.01f
C10912 XA1.XA6.MP0.G a_3440_41636# 7.76e-20
C10913 XA2.XA4.MN0.G XA2.XA1.XA5.MN0.D 0.0198f
C10914 XA6.XA3.MN0.G a_16040_44804# 0.00498f
C10915 XA0.XA9.MN1.G a_920_51140# 0.0222f
C10916 CK_SAMPLE a_16040_49732# 0.00347f
C10917 XA6.XA7.MP0.D a_16040_51844# 0.133f
C10918 XA7.XA9.MN1.G a_19928_51492# 2.84e-19
C10919 XA3.XA9.MN1.G XA5.XA1.XA5.MN2.G 4.35e-19
C10920 AVDD a_18560_49380# 0.00159f
C10921 li_9184_32484# li_9184_31872# 0.00271f
C10922 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES2.B 0.0307f
C10923 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES16.B 0.0381f
C10924 a_4808_44100# XA2.XA1.XA5.MN1.D 0.00176f
C10925 a_11000_44100# EN 0.0752f
C10926 a_17408_44100# a_18560_44100# 0.00133f
C10927 XA20.XA2a.MN0.D a_21080_42692# 0.00282f
C10928 XA20.XA3a.MN0.D XA4.XA1.XA1.MN0.S 0.0673f
C10929 XA0.XA6.MP2.G li_9184_27168# 3.5e-20
C10930 XA3.XA4.MN0.D a_8480_39876# 9.24e-20
C10931 SARN XDAC2.XC64a<0>.XRES4.B 13.9f
C10932 D<0> a_21080_50788# 0.161f
C10933 AVDD a_8480_45860# 0.00125f
C10934 XA8.XA6.MN2.D a_19928_50788# 0.0488f
C10935 a_11000_51140# XA4.XA6.MP0.G 6.76e-20
C10936 a_7328_51844# VREF 0.00396f
C10937 D<4> a_11000_50436# 0.0879f
C10938 XA4.XA6.MN2.D a_9848_50436# 0.00176f
C10939 XA0.XA6.MP2.G XA0.XA6.MN0.D 0.00148f
C10940 XDAC1.XC128a<1>.XRES16.B XDAC1.XC128a<1>.XRES1A.B 0.454f
C10941 XDAC2.XC128a<1>.XRES16.B li_14804_16728# 0.00117f
C10942 EN a_22448_41988# 5.7e-20
C10943 a_17408_43044# a_18560_43044# 0.00133f
C10944 XA0.XA6.MP0.G li_14804_6288# 0.00506f
C10945 SARN a_23600_45860# 0.0017f
C10946 VREF XA2.XA4.MN0.D 0.615f
C10947 XA20.XA3a.MN0.G a_22448_49028# 0.027f
C10948 XA0.XA4.MN0.D XA3.XA4.MN0.D 0.0342f
C10949 XA5.XA6.MP0.G a_12368_48676# 0.0881f
C10950 XA1.XA6.MP0.G a_2288_48324# 0.00417f
C10951 AVDD a_2288_43044# 0.381f
C10952 a_8480_49732# a_8480_49380# 0.0109f
C10953 a_3440_41636# a_4808_41636# 8.89e-19
C10954 SARP XDAC1.XC0.XRES8.B 27.7f
C10955 XA2.XA4.MN0.G a_4808_47620# 0.154f
C10956 VREF a_5960_46212# 0.0671f
C10957 XA0.XA7.MP0.G a_3440_43748# 0.0749f
C10958 XA2.XA1.XA5.MN2.G a_2288_43748# 0.00442f
C10959 XA8.XA1.XA5.MN2.G XA7.XA1.XA5.MP1.D 0.00329f
C10960 XA7.XA1.XA5.MN2.G XA7.XA1.XA5.MN1.D 0.0102f
C10961 AVDD a_920_40580# 0.381f
C10962 XA7.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C10963 XA8.XA12.MP0.G a_19928_53252# 0.0661f
C10964 XA0.XA12.MP0.D a_2288_52900# 0.00273f
C10965 XA0.XA12.MP0.G a_920_52900# 1.28e-19
C10966 XA5.XA11.MN1.G XA4.XA10.MP0.D 0.00744f
C10967 AVDD XA2.XA9.MN0.D 4.25e-19
C10968 a_16040_40580# a_17408_40580# 8.89e-19
C10969 XA6.XA4.MN0.G a_13520_44452# 2.2e-19
C10970 XA6.XA3.MN0.G a_14888_45860# 0.162f
C10971 XA4.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S 0.0308f
C10972 XA0.XA4.MN0.D a_920_43396# 9.14e-20
C10973 XA5.XA4.MN0.G a_14888_44452# 2.2e-19
C10974 CK_SAMPLE a_16040_50436# 0.00312f
C10975 AVDD XA8.XA6.MN0.D 3.77e-19
C10976 a_13520_52548# XA5.XA7.MP0.D 5.16e-20
C10977 a_22448_52548# a_22448_52196# 0.0109f
C10978 XA4.XA9.MN1.G a_9848_52196# 0.0862f
C10979 XB2.XA0.MP0.D CK_SAMPLE_BSSW 0.148f
C10980 XB1.XA0.MP0.D a_8408_334# 0.00524f
C10981 XB2.M1.G a_12368_n18# 0.0671f
C10982 a_12368_1390# a_13808_1390# 8e-19
C10983 XA0.XA4.MN0.D a_n232_40932# 9.25e-20
C10984 XA7.XA6.MP0.G a_12368_40228# 3.71e-19
C10985 a_n232_45156# EN 5.62e-19
C10986 XA2.XA6.MP0.G a_5960_39876# 0.00207f
C10987 XA20.XA3a.MN0.D XA8.XA1.XA4.MN0.D 1.13e-19
C10988 XA20.XA2a.MN0.D a_4808_43396# 7.39e-20
C10989 XA6.XA6.MP0.G a_16040_40228# 5.5e-19
C10990 XA2.XA4.MN0.G a_4808_41988# 1.74e-19
C10991 AVDD a_7328_46916# 0.359f
C10992 XA7.XA1.XA5.MN2.G XA6.XA6.MP2.D 0.00313f
C10993 XA6.XA9.MN1.G a_16040_50084# 0.00281f
C10994 XA1.XA9.MN1.G a_2288_49732# 0.0215f
C10995 a_22448_51140# a_23600_51140# 0.00133f
C10996 XB1.XA4.MP0.D m3_n1960_132# 0.0137f
C10997 XA20.XA2a.MN0.D a_3440_40932# 0.0733f
C10998 XA1.XA1.XA2.MP0.D a_2288_43044# 3.59e-19
C10999 XA1.XA6.MP0.G XDAC2.XC128a<1>.XRES16.B 4.21e-20
C11000 EN a_7328_42692# 0.159f
C11001 XA20.XA3a.MN0.G a_22448_50084# 0.156f
C11002 XA0.XA7.MP0.G a_920_47972# 0.00363f
C11003 D<4> a_11000_48676# 0.00918f
C11004 XA5.XA1.XA5.MN2.G XA6.XA4.MN0.G 3.9e-20
C11005 XA6.XA1.XA5.MN2.G XA5.XA4.MN0.G 0.158f
C11006 XA0.XA6.MP2.G a_920_48324# 0.0164f
C11007 XA1.XA6.MP0.G VREF 0.568f
C11008 AVDD XA8.XA1.XA5.MN1.D 0.00924f
C11009 a_8480_50084# a_9848_50084# 8.89e-19
C11010 XA0.XA6.MP0.G XA3.XA4.MN0.D 0.869f
C11011 D<0> a_21080_49028# 0.00884f
C11012 SARP SAR_IN 0.606f
C11013 D<8> XDAC2.XC128b<2>.XRES4.B 4.06e-21
C11014 a_21080_43044# XA8.XA1.XA1.MN0.S 4.06e-20
C11015 XA20.XA3.MN6.D XA8.XA3.MN0.G 0.00652f
C11016 XA1.XA6.MP0.G a_3440_46212# 7.76e-20
C11017 a_2288_48324# a_3440_48324# 0.00133f
C11018 XA5.XA1.XA5.MN2.G a_9848_44804# 1.86e-19
C11019 AVDD XA3.XA1.XA1.MN0.S 1.03f
C11020 XA1.XA4.MN0.D a_3440_47268# 0.0963f
C11021 XA8.XA4.MN0.D a_19928_47620# 0.0396f
C11022 VREF a_4808_47268# 1.19e-19
C11023 XA3.XA11.MN1.G XA4.XA11.MN1.G 0.271f
C11024 AVDD a_17408_53252# 0.361f
C11025 a_18560_53956# XA7.XA12.MP0.G 0.0688f
C11026 a_19928_53956# XA8.XA11.MN1.G 7.59e-19
C11027 XA3.XA1.XA1.MN0.S a_7328_40228# 0.0313f
C11028 XA8.XA1.XA1.MN0.S a_19928_40580# 0.00155f
C11029 XA3.XA1.XA1.MN0.D a_8480_40932# 0.0535f
C11030 a_21080_41284# a_21080_40932# 0.0109f
C11031 XA0.XA7.MP0.G a_n232_42340# 3.12e-19
C11032 XA7.XA1.XA5.MN2.G XA6.XA1.XA4.MP0.D 0.00361f
C11033 D<6> a_4808_42692# 6.49e-19
C11034 a_22448_46916# a_23600_46916# 0.00133f
C11035 AVDD a_9560_n18# 0.00236f
C11036 XA0.XA6.MP0.G a_920_43396# 5.5e-19
C11037 XA5.XA4.MN0.G a_14888_45508# 2.84e-19
C11038 XA6.XA4.MN0.G a_13520_45508# 2.84e-19
C11039 a_4808_46916# a_4808_46564# 0.0109f
C11040 a_21080_52900# a_21080_52548# 0.0109f
C11041 AVDD D<1> 2.31f
C11042 CK_SAMPLE a_11000_51140# 8.45e-19
C11043 XA8.XA10.MP0.D XA8.XA9.MN1.G 0.00406f
C11044 a_14960_3150# XB2.M1.G 2.71e-20
C11045 XB2.XA1.MN0.D XB2.XA1.MP0.D 0.208f
C11046 XB1.XA1.MN0.D a_9560_2446# 0.0727f
C11047 a_13808_2798# a_13808_2446# 0.0109f
C11048 XB1.XA1.MP0.D a_11000_2446# 3.77e-19
C11049 XB2.XA2.MN0.G XB2.XA4.MP0.D 0.0112f
C11050 SARN li_14804_32484# 0.00118f
C11051 XA0.XA6.MP0.G a_n232_40932# 3.97e-20
C11052 a_5960_45156# a_7328_45156# 8.89e-19
C11053 XA20.XA3a.MN0.D a_3440_43044# 0.0905f
C11054 XA4.XA4.MN0.G XA4.XA1.XA4.MN1.D 0.0642f
C11055 XA20.XA2a.MN0.D a_23600_44100# 0.00254f
C11056 XA1.XA4.MN0.D a_3440_41636# 9.24e-20
C11057 AVDD XA5.XA4.MN0.G 2.36f
C11058 CK_SAMPLE a_16040_48676# 6.2e-20
C11059 XA6.XA9.MN1.G a_14888_50788# 0.015f
C11060 a_3440_51492# XA2.XA1.XA5.MN2.G 0.0658f
C11061 XA3.XA7.MP0.D D<5> 2.65e-19
C11062 XA1.XA9.MN1.G a_2288_50436# 7.76e-19
C11063 XA1.XA11.MP0.D VREF 0.00176f
C11064 XDAC2.XC64b<1>.XRES16.B XDAC2.XC64b<1>.XRES1A.B 0.454f
C11065 XA0.XA6.MP2.G XDAC1.XC128a<1>.XRES16.B 0.0333f
C11066 EN XA6.XA1.XA5.MP0.D 0.0446f
C11067 a_19928_44100# XA8.XA1.XA2.MP0.D 2.92e-19
C11068 XA20.XA3a.MN0.D a_2288_40580# 0.0658f
C11069 XA20.XA2a.MN0.D a_9848_41636# 0.0144f
C11070 a_12368_43748# a_13520_43748# 0.00133f
C11071 a_n232_43748# XA0.XA1.XA5.MN0.D 0.00176f
C11072 D<4> a_9848_49732# 7.01e-19
C11073 XA0.XA6.MP2.G XA0.XA4.MN0.D 9.98f
C11074 XA7.XA1.XA5.MN2.G a_16040_49380# 0.00363f
C11075 D<0> a_21080_50084# 0.0155f
C11076 AVDD a_8480_44804# 0.00125f
C11077 li_14804_12216# li_14804_11604# 0.00271f
C11078 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES8.B 0.0228f
C11079 XDAC2.XC32a<0>.XRES16.B XDAC2.XC64a<0>.XRES16.B 0.0114f
C11080 XA0.XA4.MN0.D li_9184_6288# 0.00506f
C11081 XA0.XA1.XA4.MP1.D a_920_42340# 0.00176f
C11082 a_13520_42692# a_14888_42692# 8.89e-19
C11083 D<7> XA20.XA2a.MN0.D 0.076f
C11084 a_21080_49380# a_21080_49028# 0.0109f
C11085 XA1.XA6.MP0.G a_2288_47268# 5.95e-19
C11086 AVDD XA7.XA1.XA4.MP0.D 0.152f
C11087 XA1.XA4.MN0.D a_2288_48324# 0.0682f
C11088 XA20.XA3a.MN0.G a_23600_47972# 0.0661f
C11089 XA20.XA3.MN6.D a_22448_47972# 0.0105f
C11090 SARN a_23600_44804# 0.00206f
C11091 XA5.XA6.MP0.G a_12368_47620# 6.35e-19
C11092 D<0> XA8.XA3.MN0.G 0.534f
C11093 AVDD a_14888_53956# 0.00164f
C11094 a_12368_54308# a_13520_54308# 0.00133f
C11095 a_n232_54308# a_n232_53956# 0.0109f
C11096 SARP li_9184_22044# 0.00103f
C11097 a_n232_41284# a_920_41284# 0.00133f
C11098 XA7.XA6.MP0.G a_18560_44452# 7.76e-20
C11099 XA2.XA4.MN0.G a_5960_46564# 3.46e-19
C11100 XA8.XA4.MN0.G XA8.XA3.MN0.G 0.554f
C11101 XA8.XA7.MP0.G a_22448_43396# 0.00113f
C11102 a_16040_47620# a_16040_47268# 0.0109f
C11103 XA3.XA1.XA5.MN2.G a_4808_43044# 2.31e-19
C11104 D<4> XA4.XA1.XA2.MP0.D 0.0153f
C11105 XA3.XA6.MP0.G a_8480_44100# 7.76e-20
C11106 VREF a_7328_45156# 0.0195f
C11107 XA2.XA4.MN0.D a_4808_45156# 9.25e-20
C11108 AVDD XB2.XA2.MN0.G 0.788f
C11109 XA0.XA12.MP0.D a_3440_52196# 5.56e-19
C11110 DONE a_21080_51844# 0.0445f
C11111 XA6.XA11.MN1.G XA6.XA9.MN1.G 0.00804f
C11112 XA1.XA10.MP0.D a_2288_52900# 0.0877f
C11113 XA6.XA10.MP0.D XA7.XA10.MP0.D 0.00217f
C11114 AVDD XA7.XA8.MP0.D 0.227f
C11115 CK_SAMPLE XA4.XA7.MP0.D 0.00417f
C11116 a_9848_39876# a_11000_39876# 0.00133f
C11117 XA8.XA7.MP0.G a_21080_40932# 0.0249f
C11118 XA2.XA1.XA5.MN2.G a_4808_40580# 0.083f
C11119 SARN XB2.XA1.MN0.D 0.00249f
C11120 XA5.XA6.MP0.G a_12368_41988# 5.5e-19
C11121 XA20.XA3a.MN0.D XA8.XA1.XA5.MP1.D 0.00805f
C11122 a_11000_45860# a_11000_45508# 0.0109f
C11123 XA1.XA6.MP0.G a_2288_41636# 5.5e-19
C11124 XA2.XA4.MN0.G XA2.XA1.XA2.MP0.D 0.206f
C11125 XA6.XA3.MN0.G a_14888_44804# 0.0404f
C11126 XA7.XA9.MN1.G a_18560_51492# 0.0118f
C11127 XA3.XA9.MN1.G XA4.XA1.XA5.MN2.G 0.0494f
C11128 CK_SAMPLE a_14888_49732# 0.0693f
C11129 a_4808_51844# a_5960_51844# 0.00133f
C11130 XA6.XA7.MP0.D a_14888_51844# 0.159f
C11131 a_23600_52196# a_23600_51844# 0.0109f
C11132 a_14888_52196# XA6.XA8.MP0.D 2.11e-19
C11133 AVDD a_17408_49380# 0.356f
C11134 XA0.XA9.MN1.G a_n232_51140# 0.0469f
C11135 D<7> li_9184_27780# 0.00504f
C11136 a_4808_44804# XA2.XA1.XA2.MP0.D 2.6e-20
C11137 XA20.XA2a.MN0.D a_19928_42692# 0.00437f
C11138 XA4.XA1.XA5.MN2.D a_11000_43396# 4.58e-19
C11139 XA2.XA3.MN0.G a_4808_42340# 0.0031f
C11140 XA3.XA4.MN0.D a_7328_39876# 9.15e-20
C11141 a_9848_44100# EN 0.00576f
C11142 AVDD a_7328_45860# 0.356f
C11143 a_7328_50788# a_8480_50788# 0.00133f
C11144 a_5960_51844# VREF 0.00396f
C11145 XA0.XA6.MP2.G XA0.XA6.MP0.G 0.468f
C11146 D<4> a_9848_50436# 5.7e-19
C11147 EN a_21080_41988# 0.0739f
C11148 a_4808_43044# XA2.XA1.XA4.MN1.D 0.00176f
C11149 a_18560_49732# XA7.XA4.MN0.D 0.0659f
C11150 VREF XA1.XA4.MN0.D 0.615f
C11151 XA0.XA4.MN0.D XA2.XA4.MN0.D 0.0359f
C11152 XA0.XA6.MP2.G a_920_47268# 0.0148f
C11153 D<4> a_11000_47620# 0.0147f
C11154 AVDD a_920_43044# 0.381f
C11155 a_16040_41988# a_16040_41636# 0.0109f
C11156 VREF a_4808_46212# 7.12e-19
C11157 XA1.XA4.MN0.D a_3440_46212# 6.37e-19
C11158 XA8.XA4.MN0.D a_21080_46564# 1.28e-19
C11159 XA7.XA6.MP0.G a_18560_45508# 7.76e-20
C11160 XA4.XA6.MP0.G XA4.XA1.XA5.MN2.D 0.0325f
C11161 XA7.XA1.XA5.MN2.G XA7.XA1.XA5.MP1.D 5.21e-20
C11162 AVDD a_n232_40580# 0.00125f
C11163 a_9848_47972# a_11000_47972# 0.00133f
C11164 XA6.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C11165 XA8.XA11.MN1.G a_21080_53252# 0.0674f
C11166 XA0.XA12.MP0.D a_920_52900# 0.00183f
C11167 XA0.XA12.MP0.G a_n232_52900# 0.00258f
C11168 a_7328_53604# a_7328_53252# 0.0109f
C11169 a_17408_53604# XA7.XA11.MP0.D 0.00176f
C11170 AVDD XA2.XA9.MN1.G 0.93f
C11171 a_3440_40580# a_3440_40228# 0.0109f
C11172 a_17408_46564# a_17408_46212# 0.0109f
C11173 a_3440_46212# a_4808_46212# 8.89e-19
C11174 XA6.XA6.MP0.G XA6.XA1.XA4.MP1.D 0.00121f
C11175 XA5.XA4.MN0.G a_13520_44452# 0.00907f
C11176 XA0.XA6.MP2.G a_920_41636# 7.76e-20
C11177 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MP2.D 0.0739f
C11178 XA3.XA1.XA5.MN2.G XA4.XA1.XA1.MN0.S 5.21e-19
C11179 D<4> a_11000_41988# 7.76e-20
C11180 XA0.XA11.MN1.G a_13808_1390# 0.0021f
C11181 XA0.XA4.MN0.D a_n232_43396# 9.25e-20
C11182 VREF XA8.XA1.XA5.MP0.D 0.00202f
C11183 AVDD XA8.XA6.MP0.G 1.65f
C11184 CK_SAMPLE a_14888_50436# 0.161f
C11185 XA5.XA10.MP0.G a_13520_51844# 5.59e-19
C11186 XA4.XA9.MN1.G a_8480_52196# 2.84e-19
C11187 XB1.XA0.MP0.D CK_SAMPLE_BSSW 0.148f
C11188 XB2.XA0.MP0.D a_14960_686# 0.119f
C11189 a_8408_1390# a_8408_1038# 0.0109f
C11190 SARN XDAC2.XC128b<2>.XRES4.B 13.9f
C11191 XA20.XA2.MN1.D a_23600_44452# 0.0137f
C11192 XA8.XA1.XA5.MN2.D EN 0.122f
C11193 XA2.XA1.XA5.MN2.D XA2.XA1.XA5.MP1.D 0.0488f
C11194 XA2.XA6.MP0.G a_4808_39876# 7.76e-20
C11195 XA20.XA3a.MN0.D XA7.XA1.XA4.MN0.D 1.1e-19
C11196 XA20.XA2a.MN0.D a_3440_43396# 4.8e-20
C11197 a_23600_44804# SARP 0.066f
C11198 a_11000_44804# a_11000_44452# 0.0109f
C11199 XA6.XA6.MP0.G a_14888_40228# 7.76e-20
C11200 XA8.XA4.MN0.G a_21080_42340# 1.28e-19
C11201 XA4.XA3.MN0.G a_9848_43044# 3.62e-20
C11202 XA7.XA1.XA5.MN2.G XA6.XA6.MN2.D 6.33e-19
C11203 XA8.XA1.XA5.MN2.G D<2> 3.47e-19
C11204 a_7328_51140# XA3.XA6.MP2.D 0.00176f
C11205 XA6.XA9.MN1.G a_14888_50084# 0.00969f
C11206 a_2288_52548# VREF 0.00396f
C11207 AVDD a_5960_46916# 0.359f
C11208 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES2.B 0.0136f
C11209 XDAC1.XC128b<2>.XRES4.B XDAC1.XC128b<2>.XRES8.B 0.471f
C11210 XB1.XA4.MP0.D m3_n2104_132# 0.0273f
C11211 XA8.XA1.XA5.MN0.D XA8.XA1.XA5.MP0.D 0.00918f
C11212 XA20.XA2a.MN0.D a_2288_40932# 0.0662f
C11213 XA3.XA3.MN0.G a_9848_40580# 8.64e-19
C11214 EN a_5960_42692# 0.159f
C11215 XA4.XA6.MP0.D a_11000_49732# 0.00176f
C11216 XA1.XA6.MP0.G XA0.XA4.MN0.D 2.8e-19
C11217 XA0.XA6.MP0.D VREF 0.0115f
C11218 D<4> a_9848_48676# 3.48e-19
C11219 XA6.XA1.XA5.MN2.G XA4.XA4.MN0.G 6.95e-19
C11220 XA5.XA1.XA5.MN2.G XA5.XA4.MN0.G 0.169f
C11221 XA0.XA6.MP2.G a_n232_48324# 6.53e-19
C11222 AVDD XA7.XA1.XA5.MN1.D 0.00889f
C11223 XA0.XA6.MP0.G XA2.XA4.MN0.D 0.412f
C11224 D<0> a_19928_49028# 5.7e-19
C11225 li_9184_6900# li_9184_6288# 0.00271f
C11226 XDAC1.XC1.XRES2.B XDAC1.XC1.XRES1A.B 0.0136f
C11227 SARP XB2.XA1.MN0.D 2.94e-19
C11228 XA3.XA1.XA4.MN0.D a_8480_41988# 0.00176f
C11229 XA8.XA1.XA4.MP0.D a_21080_42340# 0.049f
C11230 a_8480_42340# a_9848_42340# 8.89e-19
C11231 XA5.XA6.MP0.G a_13520_46564# 5e-19
C11232 XA2.XA6.MP0.G XA20.XA2a.MN0.D 0.0699f
C11233 XA20.XA3a.MN0.G XA8.XA3.MN0.G 0.00217f
C11234 XA1.XA6.MP0.G a_2288_46212# 5.5e-19
C11235 a_14888_48676# a_14888_48324# 0.0109f
C11236 a_3440_48676# XA1.XA4.MN0.G 1.34e-19
C11237 XA4.XA1.XA5.MN2.G a_9848_44804# 1.95e-19
C11238 AVDD XA2.XA1.XA1.MP2.D 0.127f
C11239 XA1.XA4.MN0.D a_2288_47268# 0.0576f
C11240 VREF a_3440_47268# 1.19e-19
C11241 D<5> XA3.XA1.XA5.MN2.D 0.0285f
C11242 a_5960_53956# a_5960_53604# 0.0109f
C11243 XA3.XA11.MN1.G XA2.XA12.MP0.G 0.142f
C11244 AVDD a_16040_53252# 0.364f
C11245 a_17408_53956# XA7.XA12.MP0.G 0.0674f
C11246 a_18560_53956# XA8.XA11.MN1.G 0.0225f
C11247 SARP XDAC1.XC64a<0>.XRES4.B 13.9f
C11248 XA3.XA1.XA1.MN0.D a_7328_40932# 8.29e-20
C11249 XA7.XA1.XA5.MN2.G XA6.XA1.XA4.MN0.D 7.2e-19
C11250 XA6.XA1.XA5.MN2.G XA6.XA1.XA4.MP0.D 6.33e-19
C11251 a_13520_46916# XA5.XA3.MN0.G 0.0666f
C11252 AVDD a_8408_n18# 0.444f
C11253 XA0.XA6.MP0.G a_n232_43396# 7.76e-20
C11254 VREF a_17408_44100# 0.0251f
C11255 XA5.XA4.MN0.G a_13520_45508# 0.0104f
C11256 a_920_52548# a_2288_52548# 8.89e-19
C11257 XA4.XA10.MP0.G a_11000_52548# 0.07f
C11258 CK_SAMPLE a_9848_51140# 0.0686f
C11259 a_8480_52900# XA3.XA9.MN1.G 0.00113f
C11260 AVDD XA6.XA6.MP2.D 0.172f
C11261 a_13808_3150# XB2.M1.G 0.00116f
C11262 XB2.XA1.MN0.D SAR_IN 3.01e-19
C11263 XB1.XA1.MP0.D a_9560_2446# 0.0898f
C11264 XB1.XA1.MN0.D a_8408_2446# 0.0658f
C11265 a_8408_2798# XB1.XA4.MP0.D 0.00553f
C11266 a_9560_2798# XB1.M1.G 0.00245f
C11267 a_14960_3502# XB2.XA4.MP0.D 0.00426f
C11268 SARN li_9184_32484# 1.51e-19
C11269 D<3> a_13520_40228# 2.88e-19
C11270 XA6.XA1.XA5.MN2.D a_16040_45156# 0.155f
C11271 XA20.XA3a.MN0.D a_2288_43044# 0.00877f
C11272 D<7> a_3440_39876# 0.00173f
C11273 XA20.XA2a.MN0.D a_22448_44100# 0.00148f
C11274 XA1.XA4.MN0.D a_2288_41636# 9.15e-20
C11275 AVDD XA4.XA4.MN0.G 2.36f
C11276 CK_SAMPLE a_14888_48676# 4.46e-19
C11277 a_2288_51492# XA2.XA1.XA5.MN2.G 0.0714f
C11278 a_13520_51492# a_14888_51492# 8.89e-19
C11279 a_16040_52196# D<2> 7.56e-20
C11280 XA0.XA11.MP0.D VREF 0.00185f
C11281 EN XA6.XA1.XA5.MN0.D 0.0063f
C11282 XA1.XA6.MP0.G XDAC2.XC64b<1>.XRES16.B 4.21e-20
C11283 XA20.XA3a.MN0.D a_920_40580# 0.0674f
C11284 XA8.XA1.XA5.MN2.D a_21080_42692# 7.44e-20
C11285 XA20.XA2a.MN0.D a_8480_41636# 0.0145f
C11286 XA3.XA1.XA5.MN1.D XA3.XA1.XA5.MN0.D 0.0488f
C11287 a_n232_43748# XA0.XA1.XA2.MP0.D 0.0702f
C11288 a_22448_51140# VREF 9.95e-19
C11289 XA0.XA6.MP0.G XA1.XA6.MP0.G 6.08f
C11290 a_11000_50436# XA4.XA6.MP0.D 0.00176f
C11291 D<0> a_19928_50084# 5.7e-19
C11292 AVDD a_7328_44804# 0.356f
C11293 a_920_42692# XA0.XA1.XA4.MP0.D 0.00176f
C11294 XA5.XA1.XA4.MP1.D XA5.XA1.XA4.MP0.D 0.0488f
C11295 D<8> XDAC2.XC0.XRES4.B 0.00406f
C11296 XA0.XA6.MP2.G a_920_46212# 0.0202f
C11297 a_7328_49028# a_8480_49028# 0.00133f
C11298 AVDD XA6.XA1.XA4.MP0.D 0.152f
C11299 VREF a_2288_48324# 0.0536f
C11300 XA7.XA4.MN0.D a_18560_48676# 0.158f
C11301 XA20.XA3a.MN0.G a_22448_47972# 0.0964f
C11302 D<0> XA7.XA3.MN0.G 1.72e-19
C11303 AVDD a_13520_53956# 0.00166f
C11304 XA4.XA1.XA1.MP2.D a_11000_41284# 0.0465f
C11305 a_23600_41636# a_23600_41284# 0.0109f
C11306 XA7.XA6.MP0.G a_17408_44452# 5.5e-19
C11307 XA2.XA4.MN0.G a_4808_46564# 0.0155f
C11308 XA7.XA4.MN0.G XA8.XA3.MN0.G 0.00211f
C11309 XA8.XA4.MN0.G XA7.XA3.MN0.G 0.00211f
C11310 XA8.XA7.MP0.G a_21080_43396# 0.00442f
C11311 a_2288_47268# a_3440_47268# 0.00133f
C11312 XA2.XA1.XA5.MN2.G a_4808_43044# 0.0748f
C11313 XA3.XA6.MP0.G a_7328_44100# 5.5e-19
C11314 VREF a_5960_45156# 0.0195f
C11315 AVDD a_14960_3502# 0.468f
C11316 XA0.XA12.MP0.D a_2288_52196# 7.34e-19
C11317 DONE a_19928_51844# 0.0288f
C11318 a_13520_53252# a_13520_52900# 0.0109f
C11319 AVDD XA6.XA8.MP0.D 0.227f
C11320 CK_SAMPLE XA3.XA7.MP0.D 0.00428f
C11321 XA6.XA11.MN1.G XA5.XA9.MN0.D 1.71e-19
C11322 a_22448_40228# a_22448_39876# 0.0109f
C11323 XA8.XA1.XA5.MN2.G a_21080_40932# 1.69e-19
C11324 XA8.XA7.MP0.G a_19928_40932# 6.44e-19
C11325 XA2.XA1.XA5.MN2.G a_3440_40580# 0.00564f
C11326 XA0.XA7.MP0.G a_4808_40580# 7.1e-20
C11327 SARN SAR_IP 0.683f
C11328 XA20.XA3a.MN0.D XA8.XA1.XA5.MN1.D 0.00717f
C11329 a_22448_45860# a_23600_45860# 0.00133f
C11330 XA7.XA9.MN1.G a_17408_51492# 6.57e-19
C11331 CK_SAMPLE a_13520_49732# 0.0709f
C11332 a_12368_54308# VREF 0.00579f
C11333 AVDD a_16040_49380# 0.356f
C11334 XDAC2.XC0.XRES4.B XDAC2.XC0.XRES8.B 0.471f
C11335 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES2.B 0.0136f
C11336 XA20.XA3a.MN0.D XA3.XA1.XA1.MN0.S 0.0673f
C11337 XA0.XA6.MP2.G XDAC1.XC64b<1>.XRES16.B 3.84e-19
C11338 a_14888_45156# XA6.XA1.XA2.MP0.D 1.56e-20
C11339 XA20.XA2a.MN0.D a_18560_42692# 0.00563f
C11340 XA4.XA1.XA5.MN2.D a_9848_43396# 1.28e-19
C11341 XA2.XA3.MN0.G a_3440_42340# 4.21e-19
C11342 SARN li_14804_12216# 0.00103f
C11343 a_16040_44100# a_17408_44100# 8.89e-19
C11344 a_8480_44100# EN 0.00576f
C11345 a_3440_44100# XA1.XA1.XA5.MN1.D 0.00176f
C11346 AVDD a_5960_45860# 0.356f
C11347 XA8.XA1.XA5.MN2.G XA7.XA6.MP0.G 0.185f
C11348 XDAC2.XC128a<1>.XRES4.B XDAC2.XC32a<0>.XRES4.B 0.00284f
C11349 li_14804_17340# li_14804_16728# 0.00271f
C11350 XDAC2.XC128a<1>.XRES2.B XDAC2.XC128a<1>.XRES1A.B 0.0136f
C11351 XDAC1.XC128a<1>.XRES16.B li_9184_16728# 0.00117f
C11352 EN a_19928_41988# 1.25e-19
C11353 XA1.XA4.MN0.D XDAC1.XC128a<1>.XRES16.B 4.21e-20
C11354 XA20.XA2a.MN0.D a_14888_39876# 1.09e-19
C11355 XA3.XA1.XA2.MP0.D XA3.XA1.XA4.MN0.D 0.056f
C11356 XA7.XA1.XA2.MP0.D a_18560_42692# 0.0946f
C11357 a_16040_43044# a_17408_43044# 8.89e-19
C11358 XA0.XA6.MP0.G XDAC2.XC1.XRES16.B 0.0301f
C11359 a_17408_49732# XA7.XA4.MN0.D 0.0674f
C11360 XA0.XA4.MN0.D XA1.XA4.MN0.D 4.7f
C11361 D<0> a_21080_47972# 0.0147f
C11362 D<1> XA20.XA3a.MN0.D 0.0799f
C11363 XA0.XA6.MP2.G a_n232_47268# 3.18e-19
C11364 XA4.XA1.XA5.MN2.G a_7328_46916# 0.00455f
C11365 D<4> a_9848_47620# 5.21e-19
C11366 AVDD a_n232_43044# 0.00125f
C11367 a_7328_49732# a_7328_49380# 0.0109f
C11368 a_2288_41636# a_3440_41636# 0.00133f
C11369 a_16040_42340# XA6.XA1.XA1.MN0.S 1.34e-19
C11370 SARP li_9184_32484# 0.00103f
C11371 XA7.XA1.XA5.MN2.G XA6.XA1.XA5.MP1.D 0.00329f
C11372 XA1.XA4.MN0.G a_3440_47620# 0.154f
C11373 AVDD a_23600_40932# 0.00181f
C11374 VREF a_3440_46212# 7.12e-19
C11375 XA1.XA4.MN0.D a_2288_46212# 9.15e-20
C11376 XA8.XA4.MN0.D a_19928_46564# 4.06e-19
C11377 XA7.XA6.MP0.G a_17408_45508# 5.5e-19
C11378 XA0.XA7.MP0.G a_920_43748# 0.00442f
C11379 D<6> a_5960_44100# 7.76e-20
C11380 XA5.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C11381 XA8.XA4.MN0.G a_21080_47972# 0.155f
C11382 D<2> a_16040_44452# 1.47e-19
C11383 XA1.XA6.MP0.G a_3440_45156# 7.76e-20
C11384 XA7.XA12.MP0.G a_18560_53252# 0.0661f
C11385 XA8.XA11.MN1.G a_19928_53252# 0.0689f
C11386 AVDD XA1.XA9.MN0.D 4.25e-19
C11387 XA4.XA11.MN1.G XA4.XA10.MP0.D 0.0625f
C11388 XA3.XA12.MP0.G XA3.XA10.MP0.D 0.0632f
C11389 XA20.XA12.MP0.G a_21080_52548# 4.47e-19
C11390 XA0.XA11.MN1.G XA0.XA11.MP0.D 0.00989f
C11391 a_14888_40580# a_16040_40580# 0.00133f
C11392 XA20.XA3a.MN0.D a_8480_44804# 1.57e-20
C11393 XA6.XA6.MP0.G XA6.XA1.XA4.MN1.D 7.41e-19
C11394 XA5.XA4.MN0.G a_12368_44452# 5.54e-19
C11395 XA5.XA3.MN0.G a_13520_45860# 0.162f
C11396 XA0.XA6.MP2.G a_n232_41636# 6.49e-19
C11397 XA4.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.S 0.301f
C11398 D<4> a_9848_41988# 6.49e-19
C11399 XA0.XA11.MN1.G a_12368_1390# 0.0661f
C11400 AVDD XA7.XA6.MN0.D 3.13e-19
C11401 CK_SAMPLE a_13520_50436# 0.161f
C11402 XA8.XA9.MN1.G XA8.XA9.MN0.D 0.034f
C11403 XA3.XA9.MN1.G a_9848_52196# 2.84e-19
C11404 XA3.XA9.MN0.D a_8480_52196# 0.0492f
C11405 a_21080_52548# a_21080_52196# 0.0109f
C11406 XA5.XA10.MP0.G a_12368_51844# 0.00224f
C11407 XB2.XA0.MP0.D a_13808_686# 0.113f
C11408 XB2.XA4.MP0.D a_14960_334# 0.00258f
C11409 a_11000_1390# a_12368_1390# 8.89e-19
C11410 XA7.XA1.XA5.MN2.D EN 0.121f
C11411 XA2.XA1.XA5.MN2.D XA2.XA1.XA5.MN1.D 0.0488f
C11412 XA20.XA2.MN1.D a_22448_44452# 8.29e-20
C11413 XA20.XA3a.MN0.D XA7.XA1.XA4.MP0.D 1.1e-19
C11414 XA8.XA4.MN0.G a_19928_42340# 7.97e-19
C11415 XA1.XA4.MN0.G a_3440_41988# 1.74e-19
C11416 XA3.XA3.MN0.G a_9848_43044# 7.98e-19
C11417 a_920_52548# VREF 0.00396f
C11418 XA7.XA1.XA5.MN2.G D<2> 0.627f
C11419 a_7328_51140# D<5> 0.0688f
C11420 a_21080_51140# a_22448_51140# 8.89e-19
C11421 AVDD a_4808_46916# 0.00131f
C11422 XB1.XA4.MP0.D m3_7544_308# 0.106f
C11423 XA4.XA1.XA5.MP0.D a_11000_43396# 0.049f
C11424 XA0.XA1.XA5.MP0.D a_920_43044# 0.00176f
C11425 XA8.XA1.XA2.MP0.D XA8.XA1.XA5.MP0.D 4.34e-19
C11426 XA20.XA2a.MN0.D a_920_40932# 0.0678f
C11427 XA2.XA4.MN0.D XDAC1.XC64b<1>.XRES16.B 2.19e-20
C11428 XA3.XA3.MN0.G a_8480_40580# 0.00379f
C11429 XA8.XA6.MP0.D a_21080_50084# 0.049f
C11430 AVDD XA7.XA1.XA5.MP1.D 0.0889f
C11431 XA5.XA1.XA5.MN2.G XA4.XA4.MN0.G 0.158f
C11432 a_7328_50084# a_8480_50084# 0.00133f
C11433 XA0.XA6.MP0.G XA1.XA4.MN0.D 0.294f
C11434 D<8> li_14804_22656# 3.5e-20
C11435 SARP SAR_IP 1.01f
C11436 XA8.XA1.XA4.MP0.D a_19928_42340# 2.16e-19
C11437 XA8.XA1.XA4.MN0.D a_21080_42340# 2.16e-19
C11438 XA5.XA6.MP0.G a_12368_46564# 5.5e-19
C11439 a_920_48324# a_2288_48324# 8.89e-19
C11440 XA4.XA1.XA5.MN2.G a_8480_44804# 1.86e-19
C11441 AVDD XA2.XA1.XA1.MN0.S 1.04f
C11442 VREF a_2288_47268# 0.0191f
C11443 XA7.XA4.MN0.D a_18560_47620# 0.0396f
C11444 D<2> a_16040_45508# 0.00436f
C11445 XA1.XA12.MP0.G XA2.XA12.MP0.G 0.00217f
C11446 XA2.XA11.MN1.G XA4.XA11.MN1.G 1.54e-19
C11447 AVDD a_14888_53252# 0.00154f
C11448 a_17408_53956# XA8.XA11.MN1.G 0.0295f
C11449 a_19928_41284# a_19928_40932# 0.0109f
C11450 XA3.XA1.XA1.MP1.D a_7328_40932# 0.0465f
C11451 XA6.XA1.XA5.MN2.G XA6.XA1.XA4.MN0.D 0.00313f
C11452 a_12368_46916# XA5.XA3.MN0.G 0.0674f
C11453 a_21080_46916# a_22448_46916# 8.89e-19
C11454 XA4.XA6.MP0.G XA4.XA1.XA5.MP0.D 0.00121f
C11455 AVDD a_14960_334# 0.486f
C11456 XA20.XA3.MN6.D a_22448_43748# 5.26e-19
C11457 VREF a_16040_44100# 0.0251f
C11458 D<3> XA5.XA1.XA4.MN1.D 0.00188f
C11459 XA5.XA4.MN0.G a_12368_45508# 6.57e-19
C11460 a_3440_46916# a_3440_46564# 0.0109f
C11461 CK_SAMPLE a_8480_51140# 0.067f
C11462 XA4.XA10.MP0.G a_9848_52548# 0.128f
C11463 a_19928_52900# a_19928_52548# 0.0109f
C11464 AVDD XA6.XA6.MN2.D 3.77e-19
C11465 XB2.XA2.MN0.G XB2.M1.G 0.00145f
C11466 SAR_IP SAR_IN 0.0107f
C11467 XB1.XA1.MP0.D a_8408_2446# 0.00356f
C11468 a_12368_2798# a_12368_2446# 0.0109f
C11469 a_8408_2798# XB1.M1.G 4.74e-19
C11470 XA20.XA3a.MN0.D a_920_43044# 0.00835f
C11471 SARN XDAC2.XC0.XRES4.B 13.9f
C11472 D<3> a_12368_40228# 3.45e-20
C11473 a_23600_45508# a_23600_45156# 0.0109f
C11474 XA6.XA1.XA5.MN2.D a_14888_45156# 0.153f
C11475 a_4808_45156# a_5960_45156# 0.00133f
C11476 XA3.XA6.MP0.G XA3.XA1.XA1.MN0.D 0.00112f
C11477 XA3.XA4.MN0.G XA3.XA1.XA4.MN1.D 0.0642f
C11478 D<7> a_2288_39876# 7.77e-20
C11479 XA7.XA6.MP0.G a_18560_41284# 3.97e-20
C11480 AVDD XA3.XA4.MN0.G 2.36f
C11481 CK_SAMPLE a_13520_48676# 4.46e-19
C11482 a_920_51844# XA0.XA6.MP2.G 1.25e-19
C11483 XA0.XA11.MN1.G VREF 0.0399f
C11484 XDAC1.XC64b<1>.XRES16.B XDAC1.XC64b<1>.XRES1A.B 0.454f
C11485 XDAC2.XC64b<1>.XRES16.B li_14804_27168# 0.00117f
C11486 XA0.XA6.MP2.G li_9184_17340# 0.00508f
C11487 EN XA6.XA1.XA2.MP0.D 0.03f
C11488 XA20.XA3a.MN0.D a_n232_40580# 0.0658f
C11489 XA20.XA2a.MN0.D a_7328_41636# 0.00184f
C11490 a_11000_43748# a_12368_43748# 8.89e-19
C11491 a_21080_51140# VREF 0.00377f
C11492 XA0.XA6.MP0.G XA0.XA6.MP0.D 0.0392f
C11493 AVDD a_5960_44804# 0.356f
C11494 li_9184_12216# li_9184_11604# 0.00271f
C11495 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES8.B 0.0228f
C11496 XDAC1.XC32a<0>.XRES16.B XDAC1.XC64a<0>.XRES16.B 0.0114f
C11497 a_12368_42692# a_13520_42692# 0.00133f
C11498 XA0.XA1.XA4.MN1.D a_n232_42340# 0.00176f
C11499 XA0.XA4.MN0.D XDAC1.XC1.XRES16.B 0.0301f
C11500 D<8> XDAC1.XC0.XRES4.B 3.88e-19
C11501 D<4> a_11000_46564# 0.0695f
C11502 XA4.XA1.XA5.MN2.G a_7328_45860# 0.00363f
C11503 XA0.XA6.MP2.G a_n232_46212# 0.0141f
C11504 a_19928_49380# a_19928_49028# 0.0109f
C11505 AVDD XA6.XA1.XA4.MN0.D 0.00889f
C11506 VREF a_920_48324# 0.0536f
C11507 XA7.XA4.MN0.D a_17408_48676# 0.154f
C11508 AVDD a_12368_53956# 0.464f
C11509 a_11000_54308# a_12368_54308# 8.89e-19
C11510 XA20.XA11.MP0.D CK_SAMPLE 0.0112f
C11511 SARP XDAC1.XC128b<2>.XRES4.B 13.9f
C11512 XA4.XA1.XA1.MN0.S a_11000_41284# 0.0964f
C11513 XA1.XA4.MN0.G a_4808_46564# 2.2e-19
C11514 XA2.XA4.MN0.G a_3440_46564# 2.2e-19
C11515 XA7.XA4.MN0.G XA7.XA3.MN0.G 0.554f
C11516 XA8.XA7.MP0.G a_19928_43396# 1.95e-19
C11517 a_14888_47620# a_14888_47268# 0.0109f
C11518 XA20.XA10.MN1.D a_23600_40932# 0.00537f
C11519 XA2.XA1.XA5.MN2.G a_3440_43044# 2.31e-19
C11520 XA1.XA4.MN0.D a_3440_45156# 9.24e-20
C11521 VREF a_4808_45156# 7.39e-19
C11522 AVDD a_13808_3502# 0.00166f
C11523 XA0.XA12.MP0.D a_920_52196# 4.29e-19
C11524 XA0.XA10.MP0.D a_920_52900# 0.0893f
C11525 XA5.XA10.MP0.D XA6.XA10.MP0.D 0.00217f
C11526 AVDD XA5.XA8.MP0.D 0.227f
C11527 CK_SAMPLE XA2.XA7.MP0.D 0.00417f
C11528 XA6.XA11.MN1.G XA5.XA9.MN1.G 0.0169f
C11529 a_8480_39876# a_9848_39876# 8.89e-19
C11530 XA8.XA1.XA5.MN2.G a_19928_40932# 0.00729f
C11531 XA3.XA4.MN0.D a_8480_42692# 9.24e-20
C11532 XA2.XA1.XA5.MN2.G a_2288_40580# 0.0431f
C11533 XA0.XA7.MP0.G a_3440_40580# 0.0806f
C11534 SARN XB1.XA1.MN0.D 0.00117f
C11535 XA20.XA3a.MN0.D XA7.XA1.XA5.MN1.D 2.15e-19
C11536 a_9848_45860# a_9848_45508# 0.0109f
C11537 XA1.XA4.MN0.G XA1.XA1.XA5.MN0.D 0.0198f
C11538 XA5.XA3.MN0.G a_13520_44804# 0.0404f
C11539 a_3440_51844# a_4808_51844# 8.89e-19
C11540 XA5.XA7.MP0.D a_13520_51844# 0.159f
C11541 a_22448_52196# a_22448_51844# 0.0109f
C11542 CK_SAMPLE a_12368_49732# 0.00347f
C11543 a_11000_54308# VREF 0.00579f
C11544 a_13520_52196# XA5.XA8.MP0.D 2.11e-19
C11545 AVDD a_14888_49380# 0.00159f
C11546 XA20.XA4.MN0.D a_23600_51140# 0.0562f
C11547 D<7> XDAC1.XC64b<1>.XRES2.B 0.00405f
C11548 XA20.XA2a.MN0.D a_17408_42692# 0.00457f
C11549 XA1.XA3.MN0.G a_3440_42340# 0.0029f
C11550 XA2.XA4.MN0.D a_5960_39876# 9.14e-20
C11551 a_7328_44100# EN 0.0767f
C11552 XA3.XA6.MN2.D a_8480_50436# 0.00176f
C11553 AVDD a_4808_45860# 0.00125f
C11554 a_5960_50788# a_7328_50788# 8.89e-19
C11555 XA7.XA6.MN2.D a_18560_50788# 0.0488f
C11556 XA7.XA1.XA5.MN2.G XA7.XA6.MP0.G 0.149f
C11557 EN a_18560_41988# 1.25e-19
C11558 XA20.XA2a.MN0.D a_13520_39876# 1.09e-19
C11559 XA7.XA1.XA2.MP0.D a_17408_42692# 7.68e-20
C11560 XA3.XA1.XA2.MP0.D XA3.XA1.XA4.MP0.D 4.34e-19
C11561 a_3440_43044# XA1.XA1.XA4.MN1.D 0.00176f
C11562 D<0> a_19928_47972# 5.43e-19
C11563 XA0.XA4.MN0.D VREF 0.615f
C11564 XA3.XA1.XA5.MN2.G a_7328_46916# 7.1e-20
C11565 XA4.XA1.XA5.MN2.G a_5960_46916# 7.1e-20
C11566 AVDD a_23600_43396# 0.00154f
C11567 a_14888_41988# a_14888_41636# 0.0109f
C11568 a_2288_41988# XA1.XA1.XA1.MN0.S 3.8e-19
C11569 XA7.XA1.XA5.MN2.G XA6.XA1.XA5.MN1.D 6.68e-19
C11570 XA6.XA1.XA5.MN2.G XA6.XA1.XA5.MP1.D 5.21e-20
C11571 XA1.XA4.MN0.G a_2288_47620# 0.155f
C11572 AVDD a_22448_40932# 0.57f
C11573 VREF a_2288_46212# 0.0671f
C11574 XA3.XA4.MN0.D XA20.XA2a.MN0.D 0.073f
C11575 XA0.XA7.MP0.G a_n232_43748# 1.95e-19
C11576 a_8480_47972# a_9848_47972# 8.89e-19
C11577 D<6> a_4808_44100# 6.49e-19
C11578 XA4.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C11579 XA8.XA4.MN0.G a_19928_47972# 0.153f
C11580 D<2> a_14888_44452# 5.24e-19
C11581 XA1.XA6.MP0.G a_2288_45156# 5.5e-19
C11582 XA8.XA11.MN1.G a_18560_53252# 0.0238f
C11583 XA7.XA12.MP0.G a_17408_53252# 0.00276f
C11584 XA4.XA11.MN1.G XA3.XA10.MP0.D 0.0327f
C11585 AVDD XA1.XA9.MN1.G 0.93f
C11586 a_5960_53604# a_5960_53252# 0.0109f
C11587 a_16040_53604# XA6.XA11.MP0.D 0.00176f
C11588 a_2288_40580# a_2288_40228# 0.0109f
C11589 XA2.XA6.MP0.G a_5960_42692# 5.5e-19
C11590 a_16040_46564# a_16040_46212# 0.0109f
C11591 a_2288_46212# a_3440_46212# 0.00133f
C11592 XA5.XA3.MN0.G a_12368_45860# 0.155f
C11593 XA3.XA1.XA5.MN2.G XA3.XA1.XA1.MN0.S 0.0916f
C11594 XA0.XA11.MN1.G a_11000_1390# 0.0677f
C11595 XA20.XA3.MN0.D a_23600_43396# 0.0297f
C11596 XA3.XA9.MN1.G a_8480_52196# 0.0878f
C11597 AVDD XA7.XA6.MP0.D 0.144f
C11598 CK_SAMPLE a_12368_50436# 0.00312f
C11599 XB2.XA0.MP0.D a_12368_686# 5.79e-19
C11600 XB1.XA3.MN1.D a_9560_1038# 0.00252f
C11601 XB2.XA3.MN1.D a_14960_1390# 0.0675f
C11602 XA6.XA1.XA5.MN2.D EN 0.122f
C11603 SARN li_14804_22656# 0.00103f
C11604 XA20.XA3a.MN0.D XA6.XA1.XA4.MP0.D 1.1e-19
C11605 a_22448_44804# a_23600_44804# 0.00133f
C11606 a_9848_44804# a_9848_44452# 0.0109f
C11607 XA6.XA6.MP0.G a_12368_40228# 6.52e-20
C11608 XA1.XA4.MN0.G a_2288_41988# 5.1e-20
C11609 XA3.XA3.MN0.G a_8480_43044# 0.00291f
C11610 XA0.XA9.MN1.G a_920_49732# 0.0215f
C11611 XA6.XA1.XA5.MN2.G D<2> 0.00595f
C11612 AVDD a_3440_46916# 0.00131f
C11613 XDAC2.X16ab.XRES16.B XDAC2.XC128b<2>.XRES16.B 0.0114f
C11614 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES8.B 0.0228f
C11615 li_14804_22656# li_14804_22044# 0.00271f
C11616 XB1.XA4.MP0.D m3_7472_308# 0.0634f
C11617 XA0.XA6.MP0.G XDAC2.XC128a<1>.XRES16.B 8.44e-20
C11618 XA4.XA1.XA5.MN0.D a_11000_43396# 2.16e-19
C11619 XA4.XA1.XA5.MP0.D a_9848_43396# 2.16e-19
C11620 XA8.XA1.XA2.MP0.D XA8.XA1.XA5.MN0.D 0.056f
C11621 XA20.XA2a.MN0.D a_n232_40932# 0.0717f
C11622 XA1.XA4.MN0.D XDAC1.XC64b<1>.XRES16.B 4.21e-20
C11623 AVDD XA6.XA1.XA5.MP1.D 0.0889f
C11624 XA4.XA1.XA5.MN2.G XA4.XA4.MN0.G 0.168f
C11625 XA4.XA6.MP0.G a_11000_49732# 0.101f
C11626 XA4.XA6.MN0.D a_9848_49732# 0.00176f
C11627 XA0.XA6.MP0.G VREF 0.568f
C11628 XDAC2.XC1.XRES2.B XDAC2.XC1.XRES16.B 0.457f
C11629 XDAC2.XC1.XRES8.B XDAC2.XC1.XRES1A.B 0.0228f
C11630 EN a_n232_39876# 0.00163f
C11631 XA3.XA3.MN0.G li_14804_23076# 0.00504f
C11632 SARP XB1.XA1.MN0.D 0.00249f
C11633 XA4.XA1.XA2.MP0.D a_11000_40932# 4.25e-20
C11634 XA3.XA1.XA4.MP0.D a_7328_41988# 0.00176f
C11635 XA8.XA1.XA4.MN0.D a_19928_42340# 0.0474f
C11636 a_7328_42340# a_8480_42340# 0.00133f
C11637 a_13520_48676# a_13520_48324# 0.0109f
C11638 XA0.XA6.MP2.G a_920_45156# 6.68e-19
C11639 XA4.XA1.XA5.MN2.G a_7328_44804# 0.00486f
C11640 XA3.XA1.XA5.MN2.G a_8480_44804# 1.95e-19
C11641 AVDD XA1.XA1.XA1.MP2.D 0.127f
C11642 VREF a_920_47268# 0.0191f
C11643 XA7.XA4.MN0.D a_17408_47620# 0.00498f
C11644 D<2> a_14888_45508# 0.0031f
C11645 a_4808_53956# a_4808_53604# 0.0109f
C11646 a_18560_53956# XA7.XA11.MN1.G 0.00258f
C11647 XA2.XA11.MN1.G XA2.XA12.MP0.G 0.214f
C11648 AVDD a_13520_53252# 0.00144f
C11649 SARP li_9184_12216# 0.00103f
C11650 XA7.XA1.XA1.MN0.S a_18560_40580# 0.00155f
C11651 XA2.XA1.XA1.MN0.S a_5960_40228# 0.0313f
C11652 XA6.XA1.XA5.MN2.G XA5.XA1.XA4.MN0.D 7.72e-19
C11653 XA4.XA6.MP0.G XA4.XA1.XA5.MN0.D 7.41e-19
C11654 AVDD a_13808_334# 0.00166f
C11655 XA20.XA3a.MN0.G a_22448_43748# 0.00251f
C11656 D<3> XA5.XA1.XA4.MP1.D 7.43e-19
C11657 CK_SAMPLE a_7328_51140# 8.45e-19
C11658 XA7.XA10.MP0.D XA7.XA9.MN1.G 0.00406f
C11659 a_n232_52548# a_920_52548# 0.00133f
C11660 AVDD D<2> 2.31f
C11661 a_14960_3854# XB2.XA4.MP0.D 0.0036f
C11662 XA20.XA3a.MN0.D a_n232_43044# 0.0864f
C11663 SARN XDAC1.XC0.XRES4.B 2.01e-20
C11664 XA3.XA4.MN0.G XA3.XA1.XA4.MP1.D 0.0488f
C11665 XA2.XA3.MN0.G a_4808_43748# 0.00363f
C11666 XA7.XA6.MP0.G a_17408_41284# 4.24e-19
C11667 XA5.XA9.MN1.G a_13520_50788# 0.015f
C11668 AVDD XA2.XA4.MN0.G 2.36f
C11669 CK_SAMPLE a_12368_48676# 6.2e-20
C11670 a_920_51492# XA0.XA7.MP0.G 0.0699f
C11671 a_12368_51492# a_13520_51492# 0.00133f
C11672 XA0.XA9.MN1.G a_920_50436# 7.76e-19
C11673 EN XA5.XA1.XA5.MN0.D 0.0063f
C11674 XA20.XA2a.MN0.D a_5960_41636# 0.00184f
C11675 XA3.XA1.XA5.MN1.D XA3.XA1.XA2.MP0.D 0.0102f
C11676 XA3.XA1.XA5.MP1.D XA3.XA1.XA5.MP0.D 0.0488f
C11677 a_9848_50436# XA4.XA6.MN0.D 0.00176f
C11678 a_11000_50436# XA4.XA6.MP0.G 0.0662f
C11679 a_21080_50788# XA8.XA6.MP0.G 1.34e-19
C11680 AVDD a_4808_44804# 0.00125f
C11681 a_n232_42692# XA0.XA1.XA4.MN0.D 0.00176f
C11682 XA5.XA1.XA2.MP0.D a_13520_41636# 0.00316f
C11683 XA4.XA1.XA4.MP1.D XA4.XA1.XA4.MP0.D 0.0488f
C11684 D<8> li_14804_33096# 0.00508f
C11685 D<4> a_9848_46564# 0.0551f
C11686 XA4.XA1.XA5.MN2.G a_5960_45860# 7.1e-20
C11687 XA3.XA1.XA5.MN2.G a_7328_45860# 7.1e-20
C11688 XA0.XA6.MP2.G XA20.XA2a.MN0.D 0.0752f
C11689 a_5960_49028# a_7328_49028# 8.89e-19
C11690 AVDD XA5.XA1.XA4.MN0.D 0.00889f
C11691 D<1> XA8.XA3.MN0.G 1.72e-19
C11692 XA20.XA10.MN1.D a_23600_43396# 0.00405f
C11693 XA0.XA4.MN0.D a_920_48324# 0.0698f
C11694 AVDD a_11000_53956# 0.461f
C11695 DONE CK_SAMPLE 0.155f
C11696 XA20.XA1.MN0.D a_23600_40580# 0.0584f
C11697 XA4.XA1.XA1.MN0.S a_9848_41284# 0.0658f
C11698 a_22448_41636# a_22448_41284# 0.0109f
C11699 XA1.XA4.MN0.G a_3440_46564# 0.0155f
C11700 a_920_47268# a_2288_47268# 8.89e-19
C11701 XA8.XA1.XA5.MN2.G a_19928_43396# 0.00504f
C11702 XA20.XA10.MN1.D a_22448_40932# 1.97e-19
C11703 XA0.XA7.MP0.G a_3440_43044# 0.0732f
C11704 XA2.XA1.XA5.MN2.G a_2288_43044# 0.00551f
C11705 XA1.XA4.MN0.D a_2288_45156# 9.15e-20
C11706 VREF a_3440_45156# 7.39e-19
C11707 AVDD a_14960_3854# 0.447f
C11708 XA5.XA11.MN1.G XA5.XA9.MN0.D 1.35e-19
C11709 a_12368_53252# a_12368_52900# 0.0109f
C11710 XA0.XA10.MP0.D a_n232_52900# 0.128f
C11711 AVDD XA4.XA8.MP0.D 0.227f
C11712 CK_SAMPLE XA1.XA7.MP0.D 0.00428f
C11713 XA0.XA11.MN1.G a_n232_52548# 2.85e-19
C11714 a_n232_53604# XA0.XA9.MN1.G 7.36e-20
C11715 a_21080_40228# a_21080_39876# 0.0109f
C11716 XA8.XA1.XA5.MN2.G a_18560_40932# 0.00838f
C11717 XA3.XA4.MN0.D a_7328_42692# 9.15e-20
C11718 XA0.XA7.MP0.G a_2288_40580# 0.00417f
C11719 D<2> a_16040_41284# 7.76e-20
C11720 SARN XB1.XA1.MP0.D 0.0049f
C11721 XA20.XA3a.MN0.D XA7.XA1.XA5.MP1.D 2.15e-19
C11722 a_21080_45860# a_22448_45860# 8.89e-19
C11723 XA8.XA4.MN0.G a_21080_43748# 6.3e-19
C11724 XA1.XA4.MN0.G XA1.XA1.XA5.MP0.D 0.00138f
C11725 XA5.XA3.MN0.G a_12368_44804# 0.00498f
C11726 XA5.XA7.MP0.D a_12368_51844# 0.133f
C11727 XA2.XA9.MN1.G XA3.XA1.XA5.MN2.G 0.0494f
C11728 CK_SAMPLE a_11000_49732# 0.00347f
C11729 AVDD a_13520_49380# 0.00159f
C11730 XA20.XA4.MN0.D a_22448_51140# 3.45e-19
C11731 XDAC1.XC0.XRES4.B XDAC1.XC0.XRES8.B 0.471f
C11732 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES2.B 0.0136f
C11733 XA20.XA3a.MN0.D XA2.XA1.XA1.MN0.S 0.0673f
C11734 XA20.XA2a.MN0.D a_16040_42692# 0.00457f
C11735 XA3.XA1.XA5.MN2.D a_8480_43396# 1.28e-19
C11736 XA2.XA4.MN0.D a_4808_39876# 9.25e-20
C11737 SARN XDAC2.XC64a<0>.XRES1B.B 3.59f
C11738 a_14888_44100# a_16040_44100# 0.00133f
C11739 a_5960_44100# EN 0.0752f
C11740 a_2288_44100# XA1.XA1.XA5.MP1.D 0.00176f
C11741 XA0.XA6.MP2.G li_9184_27780# 3.5e-20
C11742 AVDD a_3440_45860# 0.00125f
C11743 XA6.XA1.XA5.MN2.G XA7.XA6.MP0.G 0.0327f
C11744 a_2288_51844# VREF 0.00396f
C11745 XDAC1.XC128a<1>.XRES4.B XDAC1.XC32a<0>.XRES4.B 0.00284f
C11746 li_9184_17340# li_9184_16728# 0.00271f
C11747 XDAC1.XC128a<1>.XRES2.B XDAC1.XC128a<1>.XRES1A.B 0.0136f
C11748 EN a_17408_41988# 0.0723f
C11749 XA0.XA4.MN0.D XDAC1.XC128a<1>.XRES16.B 8.44e-20
C11750 a_14888_43044# a_16040_43044# 0.00133f
C11751 XA0.XA6.MP0.G li_14804_6900# 0.00506f
C11752 XA0.XA6.MP0.G a_920_48324# 0.00417f
C11753 a_16040_49732# XA6.XA4.MN0.D 0.0658f
C11754 XA8.XA6.MP0.G a_21080_49028# 0.0307f
C11755 XA3.XA1.XA5.MN2.G a_5960_46916# 0.00455f
C11756 AVDD a_22448_43396# 0.438f
C11757 XA4.XA6.MP0.G a_11000_48676# 0.0881f
C11758 a_5960_49732# a_5960_49380# 0.0109f
C11759 SARP XDAC1.XC0.XRES4.B 13.9f
C11760 a_920_41636# a_2288_41636# 8.89e-19
C11761 XA2.XA3.MN0.G XDAC2.XC32a<0>.XRES1A.A 0.0138f
C11762 XA6.XA1.XA5.MN2.G XA6.XA1.XA5.MN1.D 0.0102f
C11763 AVDD a_21080_40932# 0.358f
C11764 VREF a_920_46212# 0.0671f
C11765 XA2.XA4.MN0.D XA20.XA2a.MN0.D 0.0729f
C11766 XA7.XA4.MN0.D a_18560_46564# 4.06e-19
C11767 XA3.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C11768 a_23600_53956# XA20.XA9.MP0.D 6.4e-20
C11769 CK_SAMPLE a_23600_52900# 8.74e-19
C11770 AVDD XA0.XA9.MN0.D 4.25e-19
C11771 XA7.XA11.MN1.G a_19928_53252# 2.81e-19
C11772 XA8.XA11.MN1.G a_17408_53252# 3.16e-19
C11773 a_13520_40580# a_14888_40580# 8.89e-19
C11774 XA2.XA6.MP0.G a_4808_42692# 7.76e-20
C11775 XA4.XA4.MN0.G a_11000_44452# 5.54e-19
C11776 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MP2.D 0.0736f
C11777 XA4.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S 3.84e-21
C11778 XA0.XA11.MN1.G a_9560_1390# 0.0021f
C11779 XA3.XA9.MN1.G a_7328_52196# 0.0665f
C11780 a_9848_52548# XA4.XA7.MP0.D 5.16e-20
C11781 a_19928_52548# a_19928_52196# 0.0109f
C11782 XA4.XA10.MP0.G a_11000_51844# 0.00224f
C11783 AVDD XA7.XA6.MP0.G 6.09f
C11784 CK_SAMPLE a_11000_50436# 0.00312f
C11785 XB2.M1.G a_14960_334# 3.51e-20
C11786 XB1.XA3.MN0.S a_9560_1038# 0.0288f
C11787 XB1.XA3.MN1.D a_8408_1038# 0.0114f
C11788 XB2.XA3.MN1.D a_13808_1390# 0.0535f
C11789 XB2.XA3.MN0.S a_14960_1390# 1.28e-19
C11790 a_9560_1390# a_11000_1390# 8e-19
C11791 XB1.M1.G a_11000_n18# 0.0687f
C11792 XA5.XA1.XA5.MN2.D EN 0.121f
C11793 XA8.XA1.XA5.MN2.D a_21080_44100# 0.126f
C11794 XA1.XA1.XA5.MN2.D XA1.XA1.XA5.MN1.D 0.0488f
C11795 XA20.XA3a.MN0.D XA6.XA1.XA4.MN0.D 1.1e-19
C11796 XA20.XA2a.MN0.D a_n232_43396# 7.39e-20
C11797 XA7.XA4.MN0.G a_18560_42340# 7.97e-19
C11798 XA20.XA4.MN0.D VREF 1.09e-19
C11799 XA0.XA9.MN1.G a_n232_49732# 0.00119f
C11800 XA5.XA1.XA5.MN2.G D<2> 4.48e-21
C11801 XA6.XA1.XA5.MN2.G XA5.XA6.MN2.D 6.33e-19
C11802 XA5.XA9.MN1.G a_13520_50084# 0.00969f
C11803 a_5960_51140# XA2.XA6.MP2.D 0.00176f
C11804 a_19928_51140# a_21080_51140# 0.00133f
C11805 AVDD a_2288_46916# 0.359f
C11806 XB1.XA4.MP0.D m3_n1960_1188# 0.0137f
C11807 XA4.XA1.XA5.MN0.D a_9848_43396# 0.0474f
C11808 XA0.XA1.XA5.MN0.D a_n232_43044# 0.00176f
C11809 XA0.XA1.XA2.MP0.D a_920_43044# 3.59e-19
C11810 XA20.XA2a.MN0.D XA8.XA1.XA1.MP1.D 0.0095f
C11811 EN a_2288_42692# 0.159f
C11812 AVDD XA6.XA1.XA5.MN1.D 0.00889f
C11813 XA3.XA1.XA5.MN2.G XA4.XA4.MN0.G 3.9e-20
C11814 XA4.XA1.XA5.MN2.G XA3.XA4.MN0.G 0.158f
C11815 XA8.XA7.MP0.G a_22448_48324# 8.22e-19
C11816 XA4.XA6.MP0.G a_9848_49732# 0.00239f
C11817 a_5960_50084# a_7328_50084# 8.89e-19
C11818 XA0.XA6.MP0.G XA0.XA4.MN0.D 4.81f
C11819 XA8.XA6.MP0.G a_21080_50084# 0.159f
C11820 XA8.XA6.MN0.D a_19928_50084# 0.0488f
C11821 D<8> XDAC2.XC128b<2>.XRES1B.B 4.06e-21
C11822 SARP XB1.XA1.MP0.D 0.00575f
C11823 XA1.XA6.MP0.G XA20.XA2a.MN0.D 0.0699f
C11824 a_n232_48324# a_920_48324# 0.00133f
C11825 XA0.XA6.MP2.G a_n232_45156# 7.77e-19
C11826 XA3.XA1.XA5.MN2.G a_7328_44804# 7.1e-20
C11827 XA4.XA1.XA5.MN2.G a_5960_44804# 7.1e-20
C11828 AVDD XA1.XA1.XA1.MN0.S 1.03f
C11829 XA0.XA4.MN0.D a_920_47268# 0.0576f
C11830 VREF a_n232_47268# 1.19e-19
C11831 a_17408_53956# XA7.XA11.MN1.G 0.00198f
C11832 XA2.XA11.MN1.G XA3.XA11.MN1.G 0.0251f
C11833 a_16040_53956# XA6.XA12.MP0.G 0.0658f
C11834 AVDD a_12368_53252# 0.361f
C11835 a_18560_41284# a_18560_40932# 0.0109f
C11836 XA2.XA1.XA1.MP1.D a_5960_40932# 0.0465f
C11837 XA7.XA1.XA1.MN0.S a_17408_40580# 0.0318f
C11838 XA2.XA1.XA1.MN0.S a_4808_40228# 0.0215f
C11839 XA5.XA1.XA5.MN2.G XA5.XA1.XA4.MN0.D 0.00313f
C11840 XA6.XA1.XA5.MN2.G XA5.XA1.XA4.MP0.D 0.00361f
C11841 D<7> a_3440_42692# 6.49e-19
C11842 a_11000_46916# XA4.XA3.MN0.G 0.0658f
C11843 a_19928_46916# a_21080_46916# 0.00133f
C11844 XA4.XA6.MP0.G XA4.XA1.XA2.MP0.D 0.0126f
C11845 XA4.XA4.MN0.G a_11000_45508# 6.57e-19
C11846 a_2288_46916# a_2288_46564# 0.0109f
C11847 CK_SAMPLE a_5960_51140# 8.45e-19
C11848 XA8.XA11.MN1.G XA7.XA8.MP0.D 2.37e-19
C11849 AVDD XA5.XA6.MN2.D 3.77e-19
C11850 a_18560_52900# a_18560_52548# 0.0109f
C11851 XA3.XA10.MP0.G a_8480_52548# 0.13f
C11852 a_13808_3502# XB2.M1.G 5.7e-19
C11853 a_14960_2798# XB2.XA1.MP0.D 0.0317f
C11854 a_11000_2798# a_11000_2446# 0.0109f
C11855 SARN li_14804_33096# 0.00152f
C11856 a_22448_45508# a_22448_45156# 0.0109f
C11857 XA5.XA1.XA5.MN2.D a_13520_45156# 0.153f
C11858 a_3440_45156# a_4808_45156# 8.89e-19
C11859 XA1.XA3.MN0.G a_4808_43748# 4.4e-20
C11860 XA2.XA3.MN0.G a_3440_43748# 4.21e-19
C11861 XA0.XA4.MN0.D a_920_41636# 9.14e-20
C11862 XA5.XA9.MN1.G a_12368_50788# 0.00281f
C11863 AVDD XA1.XA4.MN0.G 2.36f
C11864 CK_SAMPLE a_11000_48676# 6.2e-20
C11865 XA2.XA7.MP0.D D<6> 2.65e-19
C11866 XA0.XA9.MN1.G a_n232_50436# 0.01f
C11867 a_n232_51492# XA0.XA7.MP0.G 0.0674f
C11868 a_22448_53604# VREF 0.00125f
C11869 XDAC2.XC64b<1>.XRES4.B XDAC2.X16ab.XRES4.B 0.00284f
C11870 li_14804_27780# li_14804_27168# 0.00271f
C11871 XDAC2.XC64b<1>.XRES2.B XDAC2.XC64b<1>.XRES1A.B 0.0136f
C11872 XDAC1.XC64b<1>.XRES16.B li_9184_27168# 0.00117f
C11873 EN XA5.XA1.XA5.MP0.D 0.0446f
C11874 a_18560_44100# XA7.XA1.XA2.MP0.D 2.92e-19
C11875 XA0.XA6.MP0.G XDAC2.XC64b<1>.XRES16.B 2.4e-19
C11876 XA0.XA6.MP2.G XDAC1.XC128a<1>.XRES2.B 0.00406f
C11877 XA20.XA2a.MN0.D a_4808_41636# 0.0144f
C11878 XA3.XA1.XA5.MP1.D XA3.XA1.XA2.MP0.D 6.52e-20
C11879 a_9848_43748# a_11000_43748# 0.00133f
C11880 a_9848_50436# XA4.XA6.MP0.G 3.02e-20
C11881 D<5> a_8480_49732# 7.01e-19
C11882 a_19928_50788# XA8.XA6.MP0.G 1.75e-20
C11883 XA6.XA1.XA5.MN2.G a_12368_49380# 0.00363f
C11884 AVDD a_3440_44804# 0.00125f
C11885 XDAC2.XC64a<0>.XRES1B.B XDAC2.XC64a<0>.XRES4.B 0.428f
C11886 a_11000_42692# a_12368_42692# 8.89e-19
C11887 XA5.XA1.XA2.MP0.D a_12368_41636# 0.00224f
C11888 XA1.XA1.XA2.MP0.D XA1.XA1.XA1.MN0.S 2.11e-19
C11889 XA0.XA4.MN0.D li_9184_6900# 0.00506f
C11890 D<8> li_9184_33096# 3.45e-20
C11891 XA20.XA10.MN1.D a_22448_43396# 1.97e-19
C11892 XA3.XA1.XA5.MN2.G a_5960_45860# 0.00363f
C11893 XA6.XA4.MN0.D a_16040_48676# 0.154f
C11894 XA0.XA4.MN0.D a_n232_48324# 0.0981f
C11895 XA4.XA6.MP0.G a_11000_47620# 6.35e-19
C11896 AVDD XA5.XA1.XA4.MP0.D 0.152f
C11897 D<1> XA7.XA3.MN0.G 0.572f
C11898 XA0.XA6.MP0.G a_920_47268# 5.95e-19
C11899 a_18560_49380# a_18560_49028# 0.0109f
C11900 AVDD a_9848_53956# 0.00164f
C11901 XA20.XA11.MN0.D CK_SAMPLE 0.0826f
C11902 XA20.XA11.MP0.D a_22448_54308# 0.0467f
C11903 a_9848_54308# a_11000_54308# 0.00133f
C11904 DONE a_23600_54308# 0.0676f
C11905 SARP li_9184_22656# 0.00103f
C11906 XA8.XA1.XA1.MN0.S XA8.XA1.XA1.MP2.D 0.0708f
C11907 XA20.XA1.MN0.D a_22448_40580# 0.00246f
C11908 XA1.XA4.MN0.G a_2288_46564# 3.46e-19
C11909 XA6.XA4.MN0.G XA6.XA3.MN0.G 0.554f
C11910 a_13520_47620# a_13520_47268# 0.0109f
C11911 XA7.XA1.XA5.MN2.G a_19928_43396# 7.1e-20
C11912 XA8.XA1.XA5.MN2.G a_18560_43396# 2.66e-19
C11913 VREF a_2288_45156# 0.0195f
C11914 AVDD a_13808_3854# 0.00166f
C11915 D<5> XA3.XA1.XA5.MN0.D 0.00188f
C11916 XA5.XA11.MN1.G XA5.XA9.MN1.G 0.00349f
C11917 XA4.XA10.MP0.D XA5.XA10.MP0.D 0.00217f
C11918 AVDD XA3.XA8.MP0.D 0.227f
C11919 CK_SAMPLE XA0.XA7.MP0.D 0.00417f
C11920 a_7328_39876# a_8480_39876# 0.00133f
C11921 XA8.XA1.XA5.MN2.G a_17408_40932# 0.0245f
C11922 XA7.XA1.XA5.MN2.G a_18560_40932# 0.00631f
C11923 D<6> XA2.XA1.XA1.MN0.D 0.0192f
C11924 XA4.XA6.MP0.G a_11000_41988# 5.5e-19
C11925 XA0.XA7.MP0.G a_920_40580# 0.0506f
C11926 D<2> a_14888_41284# 6.49e-19
C11927 XA0.XA6.MP0.G a_920_41636# 5.5e-19
C11928 XA20.XA3a.MN0.D XA6.XA1.XA5.MP1.D 2.15e-19
C11929 a_8480_45860# a_8480_45508# 0.0109f
C11930 XA1.XA4.MN0.G XA1.XA1.XA2.MP0.D 0.206f
C11931 XA8.XA4.MN0.G a_19928_43748# 0.0157f
C11932 a_2288_51844# a_3440_51844# 0.00133f
C11933 a_21080_52196# a_21080_51844# 0.0109f
C11934 XA6.XA9.MN1.G a_16040_51492# 6.57e-19
C11935 CK_SAMPLE a_9848_49732# 0.0693f
C11936 XA2.XA9.MN1.G XA2.XA1.XA5.MN2.G 4.35e-19
C11937 AVDD a_12368_49380# 0.356f
C11938 a_3440_44804# XA1.XA1.XA2.MP0.D 2.6e-20
C11939 XA20.XA2a.MN0.D a_14888_42692# 0.00563f
C11940 XA3.XA1.XA5.MN2.D a_7328_43396# 4.58e-19
C11941 a_4808_44100# EN 0.00576f
C11942 D<7> li_9184_28392# 0.00504f
C11943 D<5> a_8480_50436# 5.7e-19
C11944 XA3.XA6.MP2.D a_7328_50436# 0.00176f
C11945 AVDD a_2288_45860# 0.356f
C11946 XA8.XA1.XA5.MN2.G XA6.XA6.MP0.G 3.47e-19
C11947 a_4808_50788# a_5960_50788# 0.00133f
C11948 XA7.XA6.MP2.D a_17408_50788# 0.049f
C11949 XA5.XA1.XA5.MN2.G XA7.XA6.MP0.G 0.0677f
C11950 a_920_51844# VREF 0.00396f
C11951 EN a_16040_41988# 0.0739f
C11952 a_2288_43044# XA1.XA1.XA4.MP1.D 0.00176f
C11953 XA0.XA6.MP0.G a_n232_48324# 0.00295f
C11954 a_14888_49732# XA6.XA4.MN0.D 0.0675f
C11955 a_22448_49732# VREF 0.00119f
C11956 XA8.XA6.MP0.G a_19928_49028# 0.0137f
C11957 XA8.XA7.MP0.G a_22448_47268# 6.64e-19
C11958 D<2> XA20.XA3a.MN0.D 0.0799f
C11959 AVDD a_21080_43396# 0.36f
C11960 XA4.XA6.MP0.G a_9848_48676# 0.0651f
C11961 SARP li_14804_33096# 6.57e-20
C11962 a_13520_41988# a_13520_41636# 0.0109f
C11963 XA6.XA1.XA5.MN2.G XA5.XA1.XA5.MN1.D 6.68e-19
C11964 XA0.XA4.MN0.G a_920_47620# 0.155f
C11965 AVDD a_19928_40932# 0.00154f
C11966 VREF a_n232_46212# 7.12e-19
C11967 XA0.XA4.MN0.D a_920_46212# 9.14e-20
C11968 XA1.XA4.MN0.D XA20.XA2a.MN0.D 0.073f
C11969 XA7.XA4.MN0.D a_17408_46564# 1.28e-19
C11970 a_7328_47972# a_8480_47972# 0.00133f
C11971 XA2.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C11972 XA7.XA4.MN0.G a_18560_47972# 0.153f
C11973 XA3.XA6.MP0.G XA3.XA1.XA5.MN2.D 0.0267f
C11974 a_4808_53604# a_4808_53252# 0.0109f
C11975 XA2.XA12.MP0.G XA2.XA10.MP0.D 0.0632f
C11976 XA3.XA11.MN1.G XA3.XA10.MP0.D 0.0909f
C11977 CK_SAMPLE a_22448_52900# 0.00743f
C11978 AVDD XA0.XA9.MN1.G 0.93f
C11979 XA7.XA11.MN1.G a_18560_53252# 0.0758f
C11980 a_920_40580# a_920_40228# 0.0109f
C11981 a_14888_46564# a_14888_46212# 0.0109f
C11982 a_920_46212# a_2288_46212# 8.89e-19
C11983 XA4.XA4.MN0.G a_9848_44452# 0.00907f
C11984 XA4.XA3.MN0.G a_11000_45860# 0.155f
C11985 XA8.XA7.MP0.G a_22448_41636# 9.75e-19
C11986 XA3.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S 0.327f
C11987 VREF XA7.XA1.XA5.MP0.D 0.00202f
C11988 XA4.XA10.MP0.G a_9848_51844# 5.59e-19
C11989 AVDD XA6.XA6.MP0.D 0.144f
C11990 XA7.XA9.MN1.G XA8.XA9.MN1.G 0.0531f
C11991 CK_SAMPLE a_9848_50436# 0.161f
C11992 XB1.XA3.MN0.S a_8408_1038# 0.00224f
C11993 XB2.XA3.MN0.S a_13808_1390# 0.0947f
C11994 XB1.XA0.MP0.D a_11000_686# 5.79e-19
C11995 XA4.XA1.XA5.MN2.D EN 0.122f
C11996 XA8.XA1.XA5.MN2.D a_19928_44100# 0.0877f
C11997 XA1.XA1.XA5.MN2.D XA1.XA1.XA5.MP1.D 0.0488f
C11998 SARN XDAC2.XC128b<2>.XRES1B.B 3.59f
C11999 XA5.XA6.MP0.G a_13520_40228# 3.45e-20
C12000 XA20.XA3a.MN0.D XA5.XA1.XA4.MN0.D 1.1e-19
C12001 XA20.XA2a.MN0.D XA8.XA1.XA5.MP0.D 2.15e-20
C12002 a_21080_44804# a_22448_44804# 8.89e-19
C12003 a_8480_44804# a_8480_44452# 0.0109f
C12004 XA1.XA6.MP0.G a_3440_39876# 7.76e-20
C12005 XA7.XA4.MN0.G a_17408_42340# 1.28e-19
C12006 XA0.XA4.MN0.G a_920_41988# 5.1e-20
C12007 XA8.XA10.MP0.G VREF 0.0132f
C12008 XA6.XA1.XA5.MN2.G XA5.XA6.MP2.D 0.00313f
C12009 a_21080_51492# D<0> 2.41e-19
C12010 XA5.XA9.MN1.G a_12368_50084# 0.00281f
C12011 AVDD a_920_46916# 0.359f
C12012 XDAC1.X16ab.XRES16.B XDAC1.XC128b<2>.XRES16.B 0.0114f
C12013 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES8.B 0.0228f
C12014 li_9184_22656# li_9184_22044# 0.00271f
C12015 XB1.XA4.MP0.D m3_n2104_1188# 0.0273f
C12016 XA0.XA4.MN0.D XDAC1.XC64b<1>.XRES16.B 2.4e-19
C12017 XA4.XA1.XA2.MP0.D a_9848_43396# 0.0945f
C12018 XA0.XA1.XA2.MP0.D a_n232_43044# 0.0292f
C12019 XA20.XA2a.MN0.D XA8.XA1.XA1.MN0.D 0.0224f
C12020 EN a_920_42692# 0.159f
C12021 AVDD XA5.XA1.XA5.MN1.D 0.00889f
C12022 D<1> a_18560_49028# 5.7e-19
C12023 XA4.XA1.XA5.MN2.G XA2.XA4.MN0.G 6.95e-19
C12024 XA3.XA1.XA5.MN2.G XA3.XA4.MN0.G 0.169f
C12025 XA8.XA7.MP0.G a_21080_48324# 0.00455f
C12026 D<5> a_8480_48676# 3.48e-19
C12027 a_22448_50436# VREF 0.0014f
C12028 XA8.XA6.MP0.G a_19928_50084# 6.4e-20
C12029 XDAC1.XC1.XRES2.B XDAC1.XC1.XRES16.B 0.457f
C12030 XDAC1.XC1.XRES8.B XDAC1.XC1.XRES1A.B 0.0228f
C12031 XA3.XA3.MN0.G XDAC2.X16ab.XRES1A.B 0.00405f
C12032 a_17408_43044# XA7.XA1.XA1.MN0.S 4.06e-20
C12033 XA2.XA1.XA4.MP0.D a_5960_41988# 0.00176f
C12034 XA7.XA1.XA4.MN0.D a_18560_42340# 0.0474f
C12035 a_5960_42340# a_7328_42340# 8.89e-19
C12036 a_12368_48676# a_12368_48324# 0.0109f
C12037 a_n232_48676# XA0.XA4.MN0.G 1.34e-19
C12038 D<6> XA2.XA1.XA5.MN2.D 0.0284f
C12039 XA8.XA7.MP0.G XA20.XA2.MN1.D 0.00134f
C12040 XA3.XA1.XA5.MN2.G a_5960_44804# 0.00486f
C12041 AVDD XA0.XA1.XA1.MP2.D 0.127f
C12042 XA0.XA4.MN0.D a_n232_47268# 0.0963f
C12043 XA6.XA4.MN0.D a_16040_47620# 0.00498f
C12044 XA0.XA6.MP0.G a_920_46212# 5.5e-19
C12045 a_16040_53956# XA7.XA11.MN1.G 0.0442f
C12046 a_14888_53956# XA6.XA12.MP0.G 0.0704f
C12047 XA2.XA11.MN1.G XA1.XA12.MP0.G 0.391f
C12048 AVDD a_11000_53252# 0.364f
C12049 DONE XA8.XA11.MP0.D 0.00129f
C12050 XA0.XA12.MP0.D XA2.XA12.MP0.G 0.00122f
C12051 a_3440_53956# a_3440_53604# 0.0109f
C12052 XA2.XA1.XA1.MN0.D a_5960_40932# 8.29e-20
C12053 SARP XDAC1.XC64a<0>.XRES1B.B 3.59f
C12054 XA5.XA1.XA5.MN2.G XA5.XA1.XA4.MP0.D 6.33e-19
C12055 D<7> a_2288_42692# 7.77e-20
C12056 a_9848_46916# XA4.XA3.MN0.G 0.0682f
C12057 VREF a_12368_44100# 0.0251f
C12058 XA3.XA4.MN0.D a_8480_44100# 9.24e-20
C12059 XA4.XA4.MN0.G a_9848_45508# 0.0104f
C12060 CK_SAMPLE a_4808_51140# 0.0686f
C12061 AVDD XA5.XA6.MP2.D 0.172f
C12062 XA3.XA10.MP0.G a_7328_52548# 0.0684f
C12063 a_13808_2798# XB2.XA1.MP0.D 0.0153f
C12064 XB1.XA1.MN0.D SAR_IP 3.01e-19
C12065 XA20.XA3a.MN0.D a_22448_43396# 0.0103f
C12066 SARN li_9184_33096# 4.95e-19
C12067 XA5.XA1.XA5.MN2.D a_12368_45156# 0.155f
C12068 XA2.XA4.MN0.G XA2.XA1.XA4.MP1.D 0.0488f
C12069 XA1.XA3.MN0.G a_3440_43748# 0.00371f
C12070 XA0.XA4.MN0.D a_n232_41636# 9.25e-20
C12071 AVDD XA0.XA4.MN0.G 2.36f
C12072 CK_SAMPLE a_9848_48676# 4.46e-19
C12073 a_11000_51492# a_12368_51492# 8.89e-19
C12074 a_21080_53604# VREF 0.00386f
C12075 EN XA5.XA1.XA2.MP0.D 0.03f
C12076 XA20.XA3a.MN0.D a_21080_40932# 0.0658f
C12077 XA7.XA1.XA5.MN2.D a_17408_42692# 7.44e-20
C12078 XA20.XA2a.MN0.D a_3440_41636# 0.0145f
C12079 XA8.XA1.XA5.MP1.D a_21080_43748# 0.049f
C12080 D<1> a_18560_50084# 5.7e-19
C12081 D<5> a_7328_49732# 0.0109f
C12082 XA5.XA1.XA5.MN2.G a_12368_49380# 7.1e-20
C12083 XA6.XA1.XA5.MN2.G a_11000_49380# 7.1e-20
C12084 AVDD a_2288_44804# 0.356f
C12085 a_17408_51140# VREF 0.00383f
C12086 XA4.XA1.XA4.MN1.D XA4.XA1.XA4.MN0.D 0.0488f
C12087 D<8> XDAC2.XC0.XRES1B.B 0.00406f
C12088 XA8.XA6.MP0.G a_21080_47972# 3.42e-19
C12089 XA6.XA4.MN0.D a_14888_48676# 0.158f
C12090 VREF a_22448_48676# 0.00186f
C12091 XA4.XA6.MP0.G a_9848_47620# 4.4e-19
C12092 AVDD XA4.XA1.XA4.MP0.D 0.152f
C12093 XA0.XA6.MP0.G a_n232_47268# 1.38e-19
C12094 XA7.XA6.MP0.G XA20.XA3a.MN0.D 0.0767f
C12095 a_4808_49028# a_5960_49028# 0.00133f
C12096 XA8.XA7.MP0.G a_22448_46212# 6.64e-19
C12097 AVDD a_8480_53956# 0.00166f
C12098 XA20.XA11.MN0.D a_23600_54308# 0.0852f
C12099 DONE a_22448_54308# 0.0749f
C12100 a_21080_41636# a_21080_41284# 0.0109f
C12101 XA2.XA6.MP0.G a_5960_44100# 5.5e-19
C12102 XA5.XA4.MN0.G XA6.XA3.MN0.G 0.00211f
C12103 XA6.XA4.MN0.G XA5.XA3.MN0.G 0.00211f
C12104 a_n232_47268# a_920_47268# 0.00133f
C12105 XA7.XA1.XA5.MN2.G a_18560_43396# 0.00518f
C12106 XA8.XA1.XA5.MN2.G a_17408_43396# 0.00442f
C12107 XA0.XA7.MP0.G a_920_43044# 0.00551f
C12108 XA6.XA6.MP0.G a_16040_44452# 5.5e-19
C12109 VREF a_920_45156# 0.0195f
C12110 AVDD a_9560_3150# 0.00166f
C12111 D<5> XA3.XA1.XA5.MP0.D 7.43e-19
C12112 XA4.XA12.MP0.G XA4.XA9.MN1.G 4.5e-19
C12113 a_11000_53252# a_11000_52900# 0.0109f
C12114 a_23600_53252# XA20.XA9.MP0.D 0.0341f
C12115 AVDD XA2.XA8.MP0.D 0.227f
C12116 CK_SAMPLE a_23600_52196# 7.93e-19
C12117 a_19928_40228# a_19928_39876# 0.0109f
C12118 XA7.XA1.XA5.MN2.G a_17408_40932# 0.0013f
C12119 XA2.XA4.MN0.D a_5960_42692# 9.14e-20
C12120 XA4.XA6.MP0.G a_9848_41988# 7.76e-20
C12121 XA0.XA7.MP0.G a_n232_40580# 9.86e-19
C12122 XA0.XA6.MP0.G a_n232_41636# 7.76e-20
C12123 SARN a_13808_2798# 0.00116f
C12124 XA20.XA3a.MN0.D XA6.XA1.XA5.MN1.D 2.15e-19
C12125 a_19928_45860# a_21080_45860# 0.00133f
C12126 XA4.XA3.MN0.G a_11000_44804# 0.00498f
C12127 XA4.XA7.MP0.D a_11000_51844# 0.133f
C12128 XA6.XA9.MN1.G a_14888_51492# 0.0118f
C12129 CK_SAMPLE a_8480_49732# 0.0709f
C12130 a_7328_54308# VREF 0.00579f
C12131 AVDD a_11000_49380# 0.356f
C12132 XA1.XA9.MN1.G XA3.XA1.XA5.MN2.G 4.35e-19
C12133 li_14804_33096# li_14804_32484# 0.00271f
C12134 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES8.B 0.0228f
C12135 XA20.XA3a.MN0.D XA1.XA1.XA1.MN0.S 0.0673f
C12136 XA20.XA2a.MN0.D a_13520_42692# 0.00563f
C12137 a_13520_45156# XA5.XA1.XA2.MP0.D 1.56e-20
C12138 XA1.XA4.MN0.D a_3440_39876# 9.24e-20
C12139 SARN li_14804_12636# 0.00103f
C12140 a_13520_44100# a_14888_44100# 8.89e-19
C12141 a_3440_44100# EN 0.00576f
C12142 a_920_44100# XA0.XA1.XA5.MP1.D 0.00176f
C12143 XA0.XA6.MP2.G XDAC1.XC64b<1>.XRES2.B 4.06e-21
C12144 XA7.XA1.XA5.MN2.G XA6.XA6.MP0.G 0.0959f
C12145 a_7328_51140# XA3.XA6.MP0.G 6.76e-20
C12146 D<5> a_7328_50436# 0.0863f
C12147 AVDD a_920_45860# 0.356f
C12148 D<1> a_17408_50788# 0.161f
C12149 XDAC2.XC128a<1>.XRES2.B XDAC2.XC128a<1>.XRES16.B 0.457f
C12150 XDAC2.XC128a<1>.XRES8.B XDAC2.XC128a<1>.XRES1A.B 0.0228f
C12151 EN a_14888_41988# 1.25e-19
C12152 XA20.XA2a.MN0.D a_9848_39876# 1.09e-19
C12153 a_13520_43044# a_14888_43044# 8.89e-19
C12154 XA0.XA6.MP0.G XDAC2.XC1.XRES2.B 0.00405f
C12155 a_21080_49732# VREF 0.0289f
C12156 XA8.XA7.MP0.G a_21080_47268# 0.00363f
C12157 AVDD a_19928_43396# 0.00159f
C12158 a_4808_49732# a_4808_49380# 0.0109f
C12159 D<5> a_8480_47620# 5.21e-19
C12160 SARP li_9184_33096# 0.00121f
C12161 a_n232_41636# a_920_41636# 0.00133f
C12162 a_920_41988# XA0.XA1.XA1.MN0.S 3.8e-19
C12163 XA6.XA1.XA5.MN2.G XA5.XA1.XA5.MP1.D 0.00329f
C12164 XA5.XA1.XA5.MN2.G XA5.XA1.XA5.MN1.D 0.0102f
C12165 AVDD a_18560_40932# 0.00125f
C12166 VREF XA20.XA2a.MN0.D 4.37e-19
C12167 XA0.XA4.MN0.D a_n232_46212# 6.37e-19
C12168 XA1.XA4.MN0.G XA20.XA3a.MN0.D 0.16f
C12169 XA0.XA4.MN0.G a_n232_47620# 0.154f
C12170 XA7.XA4.MN0.G a_17408_47972# 0.155f
C12171 XA6.XA6.MP0.G a_16040_45508# 5.5e-19
C12172 AVDD a_23600_52548# 0.00405f
C12173 XA3.XA11.MN1.G XA2.XA10.MP0.D 0.00744f
C12174 CK_SAMPLE a_21080_52900# 7.43e-19
C12175 a_22448_53604# a_23600_53604# 0.00133f
C12176 XA7.XA11.MN1.G a_17408_53252# 0.0762f
C12177 XA6.XA12.MP0.G a_16040_53252# 0.00276f
C12178 a_12368_40580# a_13520_40580# 0.00133f
C12179 XA20.XA3a.MN0.D a_3440_44804# 1.57e-20
C12180 XA4.XA4.MN0.G a_8480_44452# 2.2e-19
C12181 XA3.XA4.MN0.G a_9848_44452# 2.2e-19
C12182 XA4.XA3.MN0.G a_9848_45860# 0.162f
C12183 XA8.XA7.MP0.G a_21080_41636# 0.0754f
C12184 D<1> a_18560_42340# 6.49e-19
C12185 XA2.XA1.XA5.MN2.G XA2.XA1.XA1.MN0.S 0.0308f
C12186 XA0.XA11.MN1.G XB2.XA3.MN1.D 2.93e-19
C12187 D<5> a_8480_41988# 6.49e-19
C12188 XA5.XA6.MP0.G XA5.XA1.XA4.MN1.D 7.41e-19
C12189 XA20.XA3.MN6.D a_22448_43044# 7.56e-20
C12190 AVDD XA6.XA6.MN0.D 3.13e-19
C12191 XA7.XA9.MN1.G XA7.XA9.MN0.D 0.034f
C12192 a_8480_52548# XA3.XA7.MP0.D 5.16e-20
C12193 a_18560_52548# a_18560_52196# 0.0109f
C12194 CK_SAMPLE a_8480_50436# 0.161f
C12195 XB2.M1.G a_12368_334# 0.157f
C12196 a_8408_1390# a_9560_1390# 0.00133f
C12197 XB1.XA0.MP0.D a_9560_686# 0.114f
C12198 XA3.XA1.XA5.MN2.D EN 0.121f
C12199 XA5.XA6.MP0.G a_12368_40228# 2.93e-19
C12200 XA20.XA3a.MN0.D XA5.XA1.XA4.MP0.D 1.1e-19
C12201 XA20.XA2a.MN0.D XA8.XA1.XA5.MN0.D 2.15e-20
C12202 XA1.XA6.MP0.G a_2288_39876# 0.00207f
C12203 XA0.XA4.MN0.G a_n232_41988# 1.74e-19
C12204 XA7.XA10.MP0.G VREF 0.0134f
C12205 XA6.XA1.XA5.MN2.G D<3> 0.704f
C12206 XA20.XA9.MP0.D a_23600_49380# 0.00334f
C12207 a_4808_51140# XA2.XA6.MN2.D 0.00176f
C12208 a_5960_51140# D<6> 0.0672f
C12209 a_18560_51140# a_19928_51140# 8.89e-19
C12210 AVDD a_n232_46916# 0.00131f
C12211 XB1.XA4.MP0.D m3_7544_1364# 0.106f
C12212 XA20.XA2a.MN0.D XA7.XA1.XA1.MN0.D 0.022f
C12213 XA2.XA3.MN0.G a_4808_40580# 0.00359f
C12214 EN a_n232_42692# 0.0739f
C12215 AVDD XA5.XA1.XA5.MP1.D 0.0889f
C12216 D<1> a_17408_49028# 0.00884f
C12217 XA3.XA1.XA5.MN2.G XA2.XA4.MN0.G 0.158f
C12218 D<5> a_7328_48676# 0.00918f
C12219 XA3.XA6.MN0.D a_8480_49732# 0.00176f
C12220 a_4808_50084# a_5960_50084# 0.00133f
C12221 a_21080_50436# VREF 0.00393f
C12222 EN a_21080_40228# 0.0674f
C12223 D<8> li_14804_23076# 3.5e-20
C12224 XA7.XA1.XA4.MN0.D a_17408_42340# 2.16e-19
C12225 XA7.XA1.XA4.MP0.D a_18560_42340# 2.16e-19
C12226 XA3.XA1.XA5.MN2.G a_4808_44804# 1.86e-19
C12227 XA4.XA6.MP0.G a_11000_46564# 5.5e-19
C12228 AVDD XA0.XA1.XA1.MN0.S 1.04f
C12229 VREF a_22448_47620# 0.00224f
C12230 XA6.XA4.MN0.D a_14888_47620# 0.0396f
C12231 XA0.XA6.MP0.G a_n232_46212# 7.76e-20
C12232 a_14888_53956# XA7.XA11.MN1.G 0.0224f
C12233 XA0.XA12.MP0.G XA1.XA12.MP0.G 0.00217f
C12234 AVDD a_9848_53252# 0.00154f
C12235 a_17408_41284# a_17408_40932# 0.0109f
C12236 XA2.XA1.XA1.MN0.D a_4808_40932# 0.0535f
C12237 XA5.XA1.XA5.MN2.G XA4.XA1.XA4.MP0.D 0.00361f
C12238 a_18560_46916# a_19928_46916# 8.89e-19
C12239 AVDD a_9560_334# 0.00166f
C12240 VREF a_11000_44100# 0.0251f
C12241 XA3.XA4.MN0.D a_7328_44100# 9.15e-20
C12242 XA3.XA4.MN0.G a_9848_45508# 2.84e-19
C12243 XA4.XA4.MN0.G a_8480_45508# 2.84e-19
C12244 a_920_46916# a_920_46564# 0.0109f
C12245 CK_SAMPLE a_3440_51140# 0.067f
C12246 a_4808_52900# XA2.XA9.MN1.G 0.00113f
C12247 XA7.XA11.MN1.G XA7.XA8.MP0.D 6.42e-19
C12248 AVDD D<3> 2.31f
C12249 a_17408_52900# a_17408_52548# 0.0109f
C12250 XA6.XA10.MP0.D XA6.XA9.MN1.G 0.00406f
C12251 a_13808_3854# XB2.M1.G 3.5e-19
C12252 a_9560_2798# a_9560_2446# 0.0109f
C12253 XB1.XA1.MP0.D SAR_IP 0.0168f
C12254 a_14960_2798# XB2.XA1.MN0.D 0.0658f
C12255 XA20.XA3a.MN0.D a_21080_43396# 0.00756f
C12256 XA2.XA4.MN0.G XA2.XA1.XA4.MN1.D 0.0642f
C12257 a_21080_45508# a_21080_45156# 0.0109f
C12258 a_2288_45156# a_3440_45156# 0.00133f
C12259 XA0.XA6.MP2.G a_920_39876# 7.76e-20
C12260 D<4> a_11000_40228# 7.76e-20
C12261 SARN XDAC2.XC0.XRES1B.B 3.62f
C12262 AVDD a_23600_48324# 0.00181f
C12263 CK_SAMPLE a_8480_48676# 4.46e-19
C12264 XA20.XA4.MN0.D a_23600_50436# 0.00339f
C12265 XA20.XA9.MP0.D XA20.XA3.MN1.D 0.0314f
C12266 XDAC1.XC64b<1>.XRES4.B XDAC1.X16ab.XRES4.B 0.00284f
C12267 li_9184_27780# li_9184_27168# 0.00271f
C12268 XDAC1.XC64b<1>.XRES2.B XDAC1.XC64b<1>.XRES1A.B 0.0136f
C12269 XA0.XA6.MP2.G li_9184_17952# 0.00508f
C12270 XA2.XA1.XA5.MP1.D XA2.XA1.XA5.MP0.D 0.0488f
C12271 EN XA4.XA1.XA5.MP0.D 0.0446f
C12272 XA20.XA3a.MN0.D a_19928_40932# 0.0739f
C12273 XA20.XA2a.MN0.D a_2288_41636# 0.00184f
C12274 XA8.XA1.XA5.MP1.D a_19928_43748# 2.16e-19
C12275 XA8.XA1.XA5.MN1.D a_21080_43748# 2.16e-19
C12276 a_8480_43748# a_9848_43748# 8.89e-19
C12277 XA3.XA3.MN0.G XA4.XA1.XA1.MN0.S 0.00152f
C12278 a_8480_50436# XA3.XA6.MN0.D 0.00176f
C12279 XA5.XA1.XA5.MN2.G a_11000_49380# 0.00363f
C12280 AVDD a_920_44804# 0.356f
C12281 a_16040_51140# VREF 0.00383f
C12282 D<1> a_17408_50084# 0.0155f
C12283 XDAC1.XC64a<0>.XRES1B.B XDAC1.XC64a<0>.XRES4.B 0.428f
C12284 XA0.XA4.MN0.D XDAC1.XC1.XRES2.B 0.00405f
C12285 a_9848_42692# a_11000_42692# 0.00133f
C12286 D<8> XDAC1.XC0.XRES1B.B 0.0127f
C12287 XA8.XA6.MP0.G a_19928_47972# 1.28e-19
C12288 VREF a_21080_48676# 0.0188f
C12289 XA20.XA3.MN0.D a_23600_48324# 0.0836f
C12290 AVDD XA4.XA1.XA4.MN0.D 0.00889f
C12291 a_17408_49380# a_17408_49028# 0.0109f
C12292 XA8.XA7.MP0.G a_21080_46212# 0.00363f
C12293 AVDD a_7328_53956# 0.464f
C12294 XA20.XA11.MN0.D a_22448_54308# 0.00276f
C12295 DONE a_21080_54308# 0.00126f
C12296 a_23600_54660# a_23600_54308# 0.0109f
C12297 a_22448_54660# CK_SAMPLE 0.00128f
C12298 a_8480_54308# a_9848_54308# 8.89e-19
C12299 SARP XDAC1.XC128b<2>.XRES1B.B 3.59f
C12300 XA3.XA1.XA1.MP2.D a_7328_41284# 0.0465f
C12301 XA3.XA1.XA1.MN0.S a_8480_41284# 0.0674f
C12302 XA0.XA4.MN0.G a_920_46564# 3.46e-19
C12303 XA2.XA6.MP0.G a_4808_44100# 7.76e-20
C12304 XA5.XA4.MN0.G XA5.XA3.MN0.G 0.554f
C12305 a_12368_47620# a_12368_47268# 0.0109f
C12306 XA0.XA7.MP0.G a_n232_43044# 2.31e-19
C12307 XA6.XA6.MP0.G a_14888_44452# 7.76e-20
C12308 XA0.XA4.MN0.D a_920_45156# 9.14e-20
C12309 VREF a_n232_45156# 7.39e-19
C12310 AVDD a_8408_3150# 0.487f
C12311 D<5> XA3.XA1.XA2.MP0.D 0.0132f
C12312 XA20.XA10.MN1.D a_23600_52548# 0.00675f
C12313 XA5.XA11.MN1.G XA4.XA9.MN1.G 0.00116f
C12314 a_22448_53252# XA20.XA9.MP0.D 0.0215f
C12315 XA3.XA10.MP0.D XA4.XA10.MP0.D 0.00217f
C12316 AVDD XA1.XA8.MP0.D 0.227f
C12317 CK_SAMPLE a_22448_52196# 0.00664f
C12318 a_5960_39876# a_7328_39876# 8.89e-19
C12319 XA7.XA1.XA5.MN2.G a_16040_40932# 0.0256f
C12320 XA2.XA4.MN0.D a_4808_42692# 9.25e-20
C12321 SARN a_12368_2798# 0.00263f
C12322 XA20.XA3a.MN0.D XA5.XA1.XA5.MN1.D 2.15e-19
C12323 a_7328_45860# a_7328_45508# 0.0109f
C12324 XA7.XA4.MN0.G a_18560_43748# 0.0157f
C12325 XA0.XA4.MN0.G XA0.XA1.XA5.MP0.D 0.00138f
C12326 XA4.XA3.MN0.G a_9848_44804# 0.0404f
C12327 a_920_51844# a_2288_51844# 8.89e-19
C12328 XA4.XA7.MP0.D a_9848_51844# 0.159f
C12329 a_19928_52196# a_19928_51844# 0.0109f
C12330 a_9848_52196# XA4.XA8.MP0.D 2.11e-19
C12331 CK_SAMPLE a_7328_49732# 0.00347f
C12332 a_5960_54308# VREF 0.00579f
C12333 AVDD a_9848_49380# 0.00159f
C12334 XA1.XA9.MN1.G XA2.XA1.XA5.MN2.G 0.0494f
C12335 XA6.XA9.MN1.G a_13520_51492# 2.84e-19
C12336 XA20.XA2a.MN0.D a_12368_42692# 0.00457f
C12337 XA2.XA1.XA5.MN2.D a_5960_43396# 4.58e-19
C12338 D<8> a_n232_42340# 0.0031f
C12339 XA1.XA4.MN0.D a_2288_39876# 9.15e-20
C12340 SARN XDAC2.XC32a<0>.XRES1A.A 0.00394f
C12341 a_2288_44100# EN 0.0767f
C12342 D<7> XDAC1.XC64b<1>.XRES8.B 0.00687f
C12343 XA6.XA1.XA5.MN2.G XA6.XA6.MP0.G 0.00268f
C12344 AVDD a_n232_45860# 0.00125f
C12345 a_3440_50788# a_4808_50788# 8.89e-19
C12346 XA8.XA7.MP0.D VREF 0.0221f
C12347 EN a_13520_41988# 1.25e-19
C12348 XA20.XA2a.MN0.D a_8480_39876# 1.09e-19
C12349 XA6.XA1.XA2.MP0.D a_16040_42692# 7.68e-20
C12350 XA2.XA1.XA2.MP0.D XA2.XA1.XA4.MP0.D 4.34e-19
C12351 a_920_43044# XA0.XA1.XA4.MP1.D 0.00176f
C12352 a_13520_49732# XA5.XA4.MN0.D 0.0659f
C12353 a_22448_49732# a_23600_49732# 0.00133f
C12354 D<1> a_18560_47972# 5.43e-19
C12355 AVDD a_18560_43396# 0.00125f
C12356 D<5> a_7328_47620# 0.0147f
C12357 XA2.XA3.MN0.G li_14804_13248# 0.00504f
C12358 SARP XDAC2.XC0.XRES1B.B 0.00991f
C12359 a_12368_41988# a_12368_41636# 0.0109f
C12360 a_12368_42340# XA5.XA1.XA1.MN0.S 1.34e-19
C12361 XA20.XA9.MP0.D XA20.XA1.MN0.D 0.00981f
C12362 D<7> a_3440_44100# 6.49e-19
C12363 a_5960_47972# a_7328_47972# 8.89e-19
C12364 AVDD a_17408_40932# 0.358f
C12365 XA0.XA4.MN0.D XA20.XA2a.MN0.D 0.0729f
C12366 XA6.XA4.MN0.D a_16040_46564# 1.28e-19
C12367 XA0.XA6.MP0.G a_920_45156# 5.5e-19
C12368 XA0.XA4.MN0.G XA20.XA3a.MN0.D 0.138f
C12369 D<3> a_13520_44452# 5.26e-19
C12370 XA6.XA6.MP0.G a_14888_45508# 7.76e-20
C12371 XA5.XA1.XA5.MN2.G XA5.XA1.XA5.MP1.D 5.21e-20
C12372 AVDD a_22448_52548# 0.573f
C12373 a_12368_53604# XA5.XA11.MP0.D 0.00176f
C12374 a_3440_53604# a_3440_53252# 0.0109f
C12375 XA6.XA12.MP0.G a_14888_53252# 0.0661f
C12376 XA7.XA11.MN1.G a_16040_53252# 0.00648f
C12377 a_n232_40580# a_n232_40228# 0.0109f
C12378 XA3.XA4.MN0.G a_8480_44452# 0.00907f
C12379 a_13520_46564# a_13520_46212# 0.0109f
C12380 a_n232_46212# a_920_46212# 0.00133f
C12381 XA8.XA7.MP0.G a_19928_41636# 0.128f
C12382 D<1> a_17408_42340# 7.77e-20
C12383 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MP2.D 0.0739f
C12384 XA0.XA11.MN1.G XB2.XA3.MN0.S 0.00933f
C12385 XA0.XA7.MP0.G XA2.XA1.XA1.MN0.S 5.21e-19
C12386 VREF XA6.XA1.XA5.MP0.D 0.00202f
C12387 D<5> a_7328_41988# 7.77e-20
C12388 XA5.XA6.MP0.G XA5.XA1.XA4.MP1.D 0.00121f
C12389 AVDD XA6.XA6.MP0.G 5.96f
C12390 XA2.XA9.MN0.D a_4808_52196# 0.0492f
C12391 XA2.XA9.MN1.G a_5960_52196# 0.0681f
C12392 XA3.XA10.MP0.G a_8480_51844# 5.59e-19
C12393 CK_SAMPLE a_7328_50436# 0.00312f
C12394 a_14960_1742# a_14960_1390# 0.0109f
C12395 XB1.XA0.MP0.D a_8408_686# 0.118f
C12396 XB2.XA0.MP0.D a_14960_1038# 0.0794f
C12397 XA2.XA1.XA5.MN2.D EN 0.122f
C12398 XA7.XA1.XA5.MN2.D a_18560_44100# 0.0893f
C12399 XA0.XA1.XA5.MN2.D XA0.XA1.XA5.MP1.D 0.0488f
C12400 SARN li_14804_23076# 0.00103f
C12401 XA3.XA4.MN0.D XA3.XA1.XA1.MN0.D 0.00262f
C12402 XA20.XA3a.MN0.D XA4.XA1.XA4.MP0.D 1.1e-19
C12403 XA20.XA2a.MN0.D XA8.XA1.XA2.MP0.D 0.225f
C12404 a_19928_44804# a_21080_44804# 0.00133f
C12405 a_7328_44804# a_7328_44452# 0.0109f
C12406 XA1.XA6.MP0.G a_920_39876# 1.28e-19
C12407 XA6.XA4.MN0.G a_16040_42340# 1.28e-19
C12408 XA2.XA3.MN0.G a_4808_43044# 0.00321f
C12409 XA6.XA10.MP0.G VREF 0.0134f
C12410 XA5.XA1.XA5.MN2.G D<3> 0.0797f
C12411 XA20.XA10.MN1.D a_23600_48324# 0.005f
C12412 XA20.XA9.MP0.D a_22448_49380# 0.0674f
C12413 AVDD a_23600_47268# 0.00154f
C12414 XDAC2.XC128b<2>.XRES1B.B XDAC2.XC128b<2>.XRES4.B 0.428f
C12415 XB1.XA4.MP0.D m3_7472_1364# 0.0634f
C12416 a_23600_43748# a_23600_43396# 0.0109f
C12417 XA7.XA1.XA2.MP0.D XA8.XA1.XA2.MP0.D 0.00435f
C12418 XA3.XA1.XA5.MN0.D a_8480_43396# 0.0474f
C12419 XA7.XA1.XA5.MP0.D XA7.XA1.XA5.MN0.D 0.00918f
C12420 XA20.XA2a.MN0.D XA7.XA1.XA1.MP1.D 0.00946f
C12421 XA2.XA3.MN0.G a_3440_40580# 4.21e-19
C12422 EN XA8.XA1.XA4.MP1.D 0.0386f
C12423 XA2.XA1.XA5.MN2.G XA2.XA4.MN0.G 0.168f
C12424 AVDD XA4.XA1.XA5.MP1.D 0.0889f
C12425 XA7.XA6.MN0.D a_18560_50084# 0.0488f
C12426 XDAC2.XC1.XRES8.B XDAC2.XC1.XRES16.B 0.0904f
C12427 li_14804_7512# li_14804_6900# 0.00271f
C12428 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES1A.B 0.0197f
C12429 SARP a_12368_2798# 0.034f
C12430 XA2.XA1.XA4.MN0.D a_4808_41988# 0.00176f
C12431 XA7.XA1.XA4.MP0.D a_17408_42340# 0.049f
C12432 a_4808_42340# a_5960_42340# 0.00133f
C12433 D<3> a_13520_45508# 0.0031f
C12434 a_11000_48676# a_11000_48324# 0.0109f
C12435 XA8.XA7.MP0.G a_22448_45156# 8.22e-19
C12436 XA2.XA1.XA5.MN2.G a_4808_44804# 1.95e-19
C12437 XA4.XA6.MP0.G a_9848_46564# 5e-19
C12438 AVDD a_23600_41636# 0.00186f
C12439 XA20.XA3.MN0.D a_23600_47268# 0.0276f
C12440 VREF a_21080_47620# 0.067f
C12441 XA0.XA6.MP0.G XA20.XA2a.MN0.D 0.0699f
C12442 XA0.XA12.MP0.G XA2.XA11.MN1.G 1.54e-19
C12443 XA0.XA12.MP0.D XA1.XA12.MP0.G 0.278f
C12444 AVDD a_8480_53252# 0.00144f
C12445 a_2288_53956# a_2288_53604# 0.0109f
C12446 XA6.XA1.XA1.MN0.S a_16040_40580# 0.0318f
C12447 XA1.XA1.XA1.MN0.S a_3440_40228# 0.0215f
C12448 D<4> XA4.XA1.XA4.MP1.D 7.42e-19
C12449 XA3.XA4.MN0.G a_8480_45508# 0.0104f
C12450 AVDD a_8408_334# 0.487f
C12451 a_8480_46916# XA3.XA3.MN0.G 0.0666f
C12452 XA4.XA1.XA5.MN2.G XA4.XA1.XA4.MP0.D 6.33e-19
C12453 XA5.XA1.XA5.MN2.G XA4.XA1.XA4.MN0.D 7.2e-19
C12454 AVDD XA4.XA6.MP2.D 0.172f
C12455 CK_SAMPLE a_2288_51140# 8.45e-19
C12456 XA2.XA10.MP0.G a_5960_52548# 0.07f
C12457 a_12368_2798# SAR_IN 0.00271f
C12458 XB1.XA1.MP0.D XB1.XA1.MN0.D 0.208f
C12459 a_13808_2798# XB2.XA1.MN0.D 0.0974f
C12460 XA8.XA4.MN0.G a_21080_43044# 0.0222f
C12461 XA6.XA6.MP0.G a_16040_41284# 4.24e-19
C12462 XA4.XA1.XA5.MN2.D a_11000_45156# 0.155f
C12463 XA0.XA6.MP2.G a_n232_39876# 0.00197f
C12464 D<4> a_9848_40228# 6.49e-19
C12465 XA20.XA3.MN0.D a_23600_41636# 4.52e-20
C12466 SARN XDAC1.XC0.XRES1B.B 6.6e-20
C12467 XA20.XA3a.MN0.D a_19928_43396# 0.0771f
C12468 XA4.XA9.MN1.G a_11000_50788# 0.00281f
C12469 AVDD a_22448_48324# 0.416f
C12470 CK_SAMPLE a_7328_48676# 6.2e-20
C12471 XA8.XA7.MP0.D a_21080_51140# 0.00224f
C12472 a_12368_52196# D<3> 7.56e-20
C12473 a_9848_51492# a_11000_51492# 0.00133f
C12474 XA20.XA4.MN0.D a_22448_50436# 0.0215f
C12475 XA20.XA9.MP0.D XA20.XA3.MN6.D 0.343f
C12476 EN XA4.XA1.XA5.MN0.D 0.0063f
C12477 XA20.XA3a.MN0.D a_18560_40932# 0.0723f
C12478 XA6.XA1.XA5.MN2.D a_16040_42692# 7.44e-20
C12479 XA20.XA2a.MN0.D a_920_41636# 0.00184f
C12480 XA8.XA1.XA5.MN1.D a_19928_43748# 0.0494f
C12481 a_22448_50436# a_23600_50436# 0.00133f
C12482 AVDD a_n232_44804# 0.00125f
C12483 XA8.XA1.XA4.MP1.D a_21080_42692# 0.049f
C12484 XA3.XA1.XA4.MN1.D XA3.XA1.XA4.MN0.D 0.0488f
C12485 D<5> a_8480_46564# 0.0551f
C12486 VREF a_19928_48676# 1.3e-19
C12487 XA5.XA4.MN0.D a_13520_48676# 0.158f
C12488 XA20.XA3.MN0.D a_22448_48324# 0.00246f
C12489 AVDD XA3.XA1.XA4.MN0.D 0.00889f
C12490 a_3440_49028# a_4808_49028# 8.89e-19
C12491 AVDD a_5960_53956# 0.461f
C12492 XA20.XA12.MP0.G CK_SAMPLE 0.0771f
C12493 XA7.XA1.XA1.MN0.S XA8.XA1.XA1.MN0.S 0.00217f
C12494 XA3.XA1.XA1.MN0.S a_7328_41284# 0.0948f
C12495 a_19928_41636# a_19928_41284# 0.0109f
C12496 XA0.XA4.MN0.G a_n232_46564# 0.0155f
C12497 XA7.XA1.XA5.MN2.G a_16040_43396# 0.00442f
C12498 XA0.XA4.MN0.D a_n232_45156# 9.25e-20
C12499 VREF XA8.XA1.XA5.MN2.D 0.336f
C12500 AVDD XB1.XA2.MN0.G 0.788f
C12501 XA20.XA10.MN1.D a_22448_52548# 1.97e-19
C12502 a_9848_53252# a_9848_52900# 0.0109f
C12503 XA8.XA11.MP0.D a_21080_52900# 0.00176f
C12504 AVDD XA0.XA8.MP0.D 0.227f
C12505 CK_SAMPLE a_21080_52196# 0.00135f
C12506 a_18560_40228# a_18560_39876# 0.0109f
C12507 SARN a_11000_2798# 0.031f
C12508 XA20.XA3a.MN0.D XA5.XA1.XA5.MP1.D 2.15e-19
C12509 a_18560_45860# a_19928_45860# 8.89e-19
C12510 XA7.XA4.MN0.G a_17408_43748# 6.3e-19
C12511 XA0.XA4.MN0.G XA0.XA1.XA5.MN0.D 0.0198f
C12512 XA3.XA3.MN0.G a_9848_44804# 6.55e-19
C12513 XA7.XA1.XA5.MN2.G a_14888_40932# 6.44e-19
C12514 XA6.XA1.XA5.MN2.G a_16040_40932# 1.69e-19
C12515 CK_SAMPLE a_5960_49732# 0.00347f
C12516 XA5.XA9.MN1.G a_14888_51492# 2.84e-19
C12517 AVDD a_8480_49380# 0.00159f
C12518 li_9184_33096# li_9184_32484# 0.00271f
C12519 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES8.B 0.0228f
C12520 XA20.XA2a.MN0.D a_11000_42692# 0.00457f
C12521 XA2.XA1.XA5.MN2.D a_4808_43396# 1.28e-19
C12522 a_12368_44100# a_13520_44100# 0.00133f
C12523 a_920_44100# EN 0.0752f
C12524 a_n232_44100# XA0.XA1.XA5.MN1.D 0.00176f
C12525 XA0.XA6.MP2.G li_9184_28392# 3.5e-20
C12526 XA20.XA3a.MN0.D XA0.XA1.XA1.MN0.S 0.0672f
C12527 XA5.XA1.XA5.MN2.G XA6.XA6.MP0.G 1.81e-19
C12528 XA20.XA10.MN1.D a_23600_47268# 0.00423f
C12529 AVDD a_23600_46212# 0.00154f
C12530 XA20.XA9.MP0.D XA8.XA4.MN0.G 0.00237f
C12531 SARN a_23600_49380# 0.157f
C12532 XA7.XA7.MP0.D VREF 0.0234f
C12533 XA2.XA6.MP2.D a_5960_50436# 0.00176f
C12534 XA6.XA6.MP2.D a_16040_50788# 0.049f
C12535 XDAC1.XC128a<1>.XRES2.B XDAC1.XC128a<1>.XRES16.B 0.457f
C12536 XDAC1.XC128a<1>.XRES8.B XDAC1.XC128a<1>.XRES1A.B 0.0228f
C12537 EN a_12368_41988# 0.0723f
C12538 XA2.XA1.XA2.MP0.D XA2.XA1.XA4.MN0.D 0.056f
C12539 XA6.XA1.XA2.MP0.D a_14888_42692# 0.0962f
C12540 a_12368_43044# a_13520_43044# 0.00133f
C12541 XA0.XA6.MP0.G li_14804_7512# 0.00506f
C12542 a_3440_49732# a_3440_49380# 0.0109f
C12543 a_12368_49732# XA5.XA4.MN0.D 0.0674f
C12544 D<1> a_17408_47972# 0.0147f
C12545 AVDD a_17408_43396# 0.361f
C12546 XA2.XA1.XA5.MN2.G a_2288_46916# 0.00455f
C12547 D<3> XA20.XA3a.MN0.D 0.0798f
C12548 SARP XDAC1.XC0.XRES1B.B 3.6f
C12549 VREF a_22448_46564# 0.0016f
C12550 XA20.XA3.MN0.D a_23600_46212# 0.0275f
C12551 XA6.XA4.MN0.D a_14888_46564# 4.06e-19
C12552 XA20.XA10.MN1.D a_23600_41636# 0.00496f
C12553 XA0.XA6.MP0.G a_n232_45156# 7.76e-20
C12554 D<7> a_2288_44100# 7.77e-20
C12555 AVDD a_16040_40932# 0.358f
C12556 XA6.XA4.MN0.G a_16040_47972# 0.155f
C12557 D<3> a_12368_44452# 1.48e-19
C12558 XA5.XA1.XA5.MN2.G XA4.XA1.XA5.MP1.D 0.00329f
C12559 AVDD a_21080_52548# 0.405f
C12560 XA2.XA11.MN1.G XA2.XA10.MP0.D 0.0625f
C12561 XA1.XA12.MP0.G XA1.XA10.MP0.D 0.0632f
C12562 a_21080_53604# a_22448_53604# 8.89e-19
C12563 XA7.XA11.MN1.G a_14888_53252# 2.82e-19
C12564 a_11000_40580# a_12368_40580# 8.89e-19
C12565 XA3.XA3.MN0.G a_8480_45860# 0.162f
C12566 XA3.XA4.MN0.G a_7328_44452# 5.54e-19
C12567 XA1.XA6.MP0.G a_3440_42692# 7.76e-20
C12568 XA8.XA1.XA5.MN2.G a_19928_41636# 0.00417f
C12569 XA2.XA1.XA5.MN2.G XA1.XA1.XA1.MN0.S 0.301f
C12570 XA0.XA11.MN1.G XB1.XA3.MN1.D 0.00747f
C12571 XA2.XA9.MN1.G a_4808_52196# 0.0862f
C12572 AVDD XA5.XA6.MN0.D 3.13e-19
C12573 a_17408_52548# a_17408_52196# 0.0109f
C12574 XA3.XA10.MP0.G a_7328_51844# 0.00224f
C12575 CK_SAMPLE a_5960_50436# 0.00312f
C12576 XB2.XA4.MP0.D CK_SAMPLE_BSSW 0.00524f
C12577 XB2.XA0.MP0.D a_13808_1038# 0.158f
C12578 XA20.XA3a.MN0.D XA4.XA1.XA4.MN0.D 1.1e-19
C12579 XA6.XA4.MN0.G a_14888_42340# 7.97e-19
C12580 XA1.XA3.MN0.G a_4808_43044# 4.4e-20
C12581 XA2.XA3.MN0.G a_3440_43044# 4.21e-19
C12582 XA0.XA1.XA5.MN2.D XA0.XA1.XA5.MN1.D 0.0488f
C12583 XA7.XA1.XA5.MN2.D a_17408_44100# 0.124f
C12584 XA1.XA1.XA5.MN2.D EN 0.121f
C12585 XA20.XA10.MN1.D a_22448_48324# 1.78e-19
C12586 XA4.XA9.MN1.G a_11000_50084# 0.00281f
C12587 SARN XA20.XA3.MN1.D 0.143f
C12588 a_17408_51140# a_18560_51140# 0.00133f
C12589 XA5.XA1.XA5.MN2.G XA4.XA6.MP2.D 0.00313f
C12590 AVDD a_22448_47268# 0.404f
C12591 XA5.XA10.MP0.G VREF 0.0134f
C12592 XB1.XA4.MP0.D m3_n1960_2244# 0.0137f
C12593 XA1.XA3.MN0.G a_3440_40580# 0.00379f
C12594 XA3.XA1.XA5.MP0.D a_8480_43396# 2.16e-19
C12595 XA3.XA1.XA5.MN0.D a_7328_43396# 2.16e-19
C12596 XA7.XA1.XA2.MP0.D XA7.XA1.XA5.MN0.D 0.056f
C12597 XA20.XA2a.MN0.D XA6.XA1.XA1.MP1.D 0.00946f
C12598 EN XA8.XA1.XA4.MN1.D 3.17e-19
C12599 XA3.XA6.MP0.G a_8480_49732# 0.00239f
C12600 XA3.XA6.MP0.D a_7328_49732# 0.00176f
C12601 XA0.XA7.MP0.G XA2.XA4.MN0.G 3.9e-20
C12602 XA2.XA1.XA5.MN2.G XA1.XA4.MN0.G 0.158f
C12603 AVDD XA4.XA1.XA5.MN1.D 0.00889f
C12604 a_3440_50084# a_4808_50084# 8.89e-19
C12605 D<8> XDAC2.X16ab.XRES1A.B 4.06e-21
C12606 SARP a_11000_2798# 0.00529f
C12607 a_16040_43044# XA6.XA1.XA1.MN0.S 4.06e-20
C12608 D<3> a_12368_45508# 0.00436f
C12609 a_22448_48676# a_23600_48676# 0.00133f
C12610 XA8.XA7.MP0.G a_21080_45156# 0.00486f
C12611 XA2.XA1.XA5.MN2.G a_3440_44804# 1.86e-19
C12612 AVDD a_22448_41636# 0.569f
C12613 XA7.XA6.MP0.G XA7.XA3.MN0.G 0.05f
C12614 XA5.XA4.MN0.D a_13520_47620# 0.0396f
C12615 VREF a_19928_47620# 7.12e-19
C12616 XA0.XA12.MP0.D XA2.XA11.MN1.G 0.271f
C12617 a_14888_53956# XA6.XA11.MN1.G 7.59e-19
C12618 a_13520_53956# XA5.XA12.MP0.G 0.0688f
C12619 AVDD a_7328_53252# 0.361f
C12620 a_16040_41284# a_16040_40932# 0.0109f
C12621 XA1.XA1.XA1.MN0.D a_3440_40932# 0.0535f
C12622 XA6.XA1.XA1.MN0.S a_14888_40580# 0.00155f
C12623 XA1.XA1.XA1.MN0.S a_2288_40228# 0.0313f
C12624 SARP XDAC1.XC32a<0>.XRES1A.A 0.00394f
C12625 XA2.XA4.MN0.D a_5960_44100# 9.14e-20
C12626 XA3.XA6.MP0.G XA3.XA1.XA5.MN0.D 7.41e-19
C12627 XA3.XA4.MN0.G a_7328_45508# 6.57e-19
C12628 a_n232_46916# a_n232_46564# 0.0109f
C12629 AVDD CK_SAMPLE_BSSW 14.7f
C12630 a_17408_46916# a_18560_46916# 0.00133f
C12631 a_7328_46916# XA3.XA3.MN0.G 0.0674f
C12632 XA4.XA1.XA5.MN2.G XA4.XA1.XA4.MN0.D 0.00313f
C12633 D<4> XA4.XA1.XA4.MN1.D 0.00188f
C12634 a_16040_52900# a_16040_52548# 0.0109f
C12635 XA2.XA10.MP0.G a_4808_52548# 0.128f
C12636 CK_SAMPLE a_920_51140# 8.45e-19
C12637 AVDD XA4.XA6.MN2.D 3.77e-19
C12638 a_8408_2798# a_8408_2446# 0.0109f
C12639 XA8.XA4.MN0.G a_19928_43044# 0.0409f
C12640 XA1.XA4.MN0.G XA1.XA1.XA4.MN1.D 0.0642f
C12641 XA6.XA6.MP0.G a_14888_41284# 3.97e-20
C12642 a_19928_45508# a_19928_45156# 0.0109f
C12643 XA4.XA1.XA5.MN2.D a_9848_45156# 0.153f
C12644 a_920_45156# a_2288_45156# 8.89e-19
C12645 XA2.XA6.MP0.G XA2.XA1.XA1.MN0.D 0.00159f
C12646 XA20.XA3a.MN0.D a_18560_43396# 0.0723f
C12647 XA4.XA9.MN1.G a_9848_50788# 0.015f
C12648 CK_SAMPLE a_5960_48676# 6.2e-20
C12649 AVDD a_21080_48324# 0.359f
C12650 XA8.XA7.MP0.D a_19928_51140# 0.00388f
C12651 XA1.XA7.MP0.D D<7> 2.65e-19
C12652 a_17408_53604# VREF 0.00396f
C12653 XA20.XA9.MP0.D XA20.XA3a.MN0.G 0.519f
C12654 XDAC2.XC64b<1>.XRES8.B XDAC2.XC64b<1>.XRES1A.B 0.0228f
C12655 XDAC2.XC64b<1>.XRES2.B XDAC2.XC64b<1>.XRES16.B 0.457f
C12656 XA0.XA6.MP2.G XDAC1.XC128a<1>.XRES8.B 0.00688f
C12657 EN XA4.XA1.XA2.MP0.D 0.03f
C12658 XA2.XA1.XA5.MN1.D XA2.XA1.XA5.MN0.D 0.0488f
C12659 XA2.XA1.XA5.MP1.D XA2.XA1.XA2.MP0.D 6.52e-20
C12660 XA20.XA3a.MN0.D a_17408_40932# 0.0674f
C12661 XA20.XA2a.MN0.D a_n232_41636# 0.0144f
C12662 a_7328_43748# a_8480_43748# 0.00133f
C12663 XA3.XA3.MN0.G XA3.XA1.XA1.MN0.S 0.00995f
C12664 XA20.XA10.MN1.D a_23600_46212# 0.00423f
C12665 AVDD XA20.XA2.MN1.D 0.461f
C12666 a_8480_50436# XA3.XA6.MP0.G 3.02e-20
C12667 a_7328_50436# XA3.XA6.MP0.D 0.00176f
C12668 a_18560_50788# XA7.XA6.MP0.G 1.75e-20
C12669 li_14804_12636# li_14804_12216# 0.00411f
C12670 XDAC2.XC32a<0>.XRES2.B XDAC2.XC64a<0>.XRES2.B 1.67e-19
C12671 XA0.XA4.MN0.D li_9184_7512# 0.00506f
C12672 a_8480_42692# a_9848_42692# 8.89e-19
C12673 XA8.XA1.XA2.MP0.D a_21080_41988# 0.0219f
C12674 XA4.XA1.XA2.MP0.D a_11000_41636# 0.00224f
C12675 XA8.XA1.XA4.MN1.D a_21080_42692# 2.16e-19
C12676 XA8.XA1.XA4.MP1.D a_19928_42692# 2.16e-19
C12677 XA2.XA1.XA5.MN2.G a_2288_45860# 0.00363f
C12678 D<5> a_7328_46564# 0.0695f
C12679 VREF a_18560_48676# 1.3e-19
C12680 XA5.XA4.MN0.D a_12368_48676# 0.154f
C12681 AVDD XA3.XA1.XA4.MP0.D 0.152f
C12682 D<1> XA3.XA3.MN0.G 0.0363f
C12683 D<2> XA6.XA3.MN0.G 0.572f
C12684 XA6.XA6.MP0.G XA20.XA3a.MN0.D 0.0771f
C12685 a_16040_49380# a_16040_49028# 0.0109f
C12686 AVDD a_4808_53956# 0.00164f
C12687 XA20.XA12.MP0.D CK_SAMPLE 0.155f
C12688 a_22448_54660# a_22448_54308# 0.0109f
C12689 XA20.XA12.MP0.G a_23600_54308# 2.99e-19
C12690 a_7328_54308# a_8480_54308# 0.00133f
C12691 SARP li_9184_23076# 0.00103f
C12692 XA7.XA1.XA1.MN0.S XA7.XA1.XA1.MP2.D 0.0708f
C12693 XA20.XA3a.MN0.D a_23600_47268# 0.0158f
C12694 XA4.XA4.MN0.G XA4.XA3.MN0.G 0.554f
C12695 a_11000_47620# a_11000_47268# 0.0109f
C12696 XA7.XA1.XA5.MN2.G a_14888_43396# 1.95e-19
C12697 D<1> a_18560_43748# 6.49e-19
C12698 VREF XA7.XA1.XA5.MN2.D 0.341f
C12699 XA20.XA3.MN0.D XA20.XA2.MN1.D 0.617f
C12700 AVDD a_9560_3502# 0.00166f
C12701 SARN XA20.XA1.MN0.D 3.99e-19
C12702 XA4.XA11.MN1.G XA4.XA9.MN1.G 0.00804f
C12703 a_21080_53252# XA8.XA10.MP0.D 0.0661f
C12704 XA2.XA10.MP0.D XA3.XA10.MP0.D 0.00217f
C12705 AVDD a_23600_51844# 0.00186f
C12706 CK_SAMPLE a_19928_52196# 6.74e-19
C12707 a_4808_39876# a_5960_39876# 0.00133f
C12708 XA1.XA4.MN0.D a_3440_42692# 9.24e-20
C12709 XA20.XA3a.MN0.D XA4.XA1.XA5.MP1.D 2.15e-19
C12710 a_5960_45860# a_5960_45508# 0.0109f
C12711 D<3> a_13520_41284# 6.49e-19
C12712 XA0.XA4.MN0.G XA0.XA1.XA2.MP0.D 0.206f
C12713 XA3.XA3.MN0.G a_8480_44804# 0.0433f
C12714 D<7> XA1.XA1.XA1.MN0.D 0.0166f
C12715 XA6.XA1.XA5.MN2.G a_14888_40932# 0.00729f
C12716 a_8480_52196# XA3.XA8.MP0.D 2.11e-19
C12717 CK_SAMPLE a_4808_49732# 0.0693f
C12718 XA5.XA9.MN1.G a_13520_51492# 0.0118f
C12719 AVDD a_7328_49380# 0.356f
C12720 a_17408_52548# XA8.XA1.XA5.MN2.G 1.75e-19
C12721 a_18560_52196# a_18560_51844# 0.0109f
C12722 XA3.XA7.MP0.D a_8480_51844# 0.159f
C12723 a_n232_51844# a_920_51844# 0.00133f
C12724 XA20.XA2a.MN0.D a_9848_42692# 0.00563f
C12725 XA8.XA1.XA5.MN2.D XA8.XA1.XA2.MP0.D 4.72e-19
C12726 D<7> li_9184_29004# 0.00504f
C12727 a_n232_44100# EN 0.0767f
C12728 a_2288_50788# a_3440_50788# 0.00133f
C12729 XA20.XA10.MN1.D a_22448_47268# 2.14e-19
C12730 AVDD a_22448_46212# 0.368f
C12731 XA6.XA7.MP0.D VREF 0.0234f
C12732 a_21080_51492# XA8.XA6.MP0.G 4.06e-20
C12733 a_n232_43044# XA0.XA1.XA4.MN1.D 0.00176f
C12734 EN a_11000_41988# 0.0739f
C12735 a_17408_49732# VREF 0.029f
C12736 a_21080_49732# a_22448_49732# 8.89e-19
C12737 XA3.XA6.MP0.G a_8480_48676# 0.0651f
C12738 AVDD a_16040_43396# 0.361f
C12739 XA0.XA7.MP0.G a_2288_46916# 7.1e-20
C12740 XA2.XA1.XA5.MN2.G a_920_46916# 7.1e-20
C12741 XA7.XA6.MP0.G a_18560_49028# 0.0137f
C12742 XA2.XA3.MN0.G XDAC2.XC32a<0>.XRES16.B 0.0186f
C12743 a_11000_41988# a_11000_41636# 0.0109f
C12744 VREF a_21080_46564# 0.0171f
C12745 XA20.XA10.MN1.D a_22448_41636# 1.97e-19
C12746 a_4808_47972# a_5960_47972# 0.00133f
C12747 AVDD a_14888_40932# 0.00125f
C12748 XA2.XA6.MP0.G XA2.XA1.XA5.MN2.D 0.0268f
C12749 XA6.XA4.MN0.G a_14888_47972# 0.153f
C12750 a_23600_48324# a_23600_47972# 0.0109f
C12751 a_22448_48324# XA20.XA3a.MN0.D 9.13e-20
C12752 XA4.XA1.XA5.MN2.G XA4.XA1.XA5.MP1.D 5.21e-20
C12753 XA5.XA1.XA5.MN2.G XA4.XA1.XA5.MN1.D 6.68e-19
C12754 AVDD a_19928_52548# 0.00166f
C12755 a_11000_53604# XA4.XA11.MP0.D 0.00176f
C12756 a_2288_53604# a_2288_53252# 0.0109f
C12757 XA2.XA11.MN1.G XA1.XA10.MP0.D 0.0327f
C12758 XA6.XA11.MN1.G a_16040_53252# 0.0674f
C12759 a_23600_40932# a_23600_40580# 0.0109f
C12760 a_12368_46564# a_12368_46212# 0.0109f
C12761 XA3.XA3.MN0.G a_7328_45860# 0.155f
C12762 XA1.XA6.MP0.G a_2288_42692# 5.5e-19
C12763 XA8.XA1.XA5.MN2.G a_18560_41636# 0.131f
C12764 XA0.XA11.MN1.G XB1.XA3.MN0.S 0.00933f
C12765 XA0.XA7.MP0.G XA1.XA1.XA1.MN0.S 0.0916f
C12766 XA2.XA9.MN1.G a_3440_52196# 2.84e-19
C12767 XA6.XA9.MN1.G XA7.XA9.MN1.G 0.00217f
C12768 CK_SAMPLE a_4808_50436# 0.161f
C12769 AVDD XA5.XA6.MP0.D 0.144f
C12770 XB2.XA4.MP0.D a_14960_686# 0.0023f
C12771 XB1.XA3.MN1.D a_9560_1390# 0.0535f
C12772 a_13808_1742# a_13808_1390# 0.0109f
C12773 SARN XDAC2.X16ab.XRES1A.B 3.59f
C12774 XA0.XA6.MP0.G a_2288_39876# 1.28e-19
C12775 XA20.XA3a.MN0.D XA3.XA1.XA4.MN0.D 1.1e-19
C12776 a_18560_44804# a_19928_44804# 8.89e-19
C12777 a_5960_44804# a_5960_44452# 0.0109f
C12778 XA8.XA3.MN0.G a_19928_43396# 6.8e-20
C12779 XA1.XA3.MN0.G a_3440_43044# 0.00291f
C12780 XA0.XA1.XA5.MN2.D EN 0.162f
C12781 XA4.XA9.MN1.G a_9848_50084# 0.00969f
C12782 SARN XA20.XA3.MN6.D 0.0502f
C12783 a_3440_51140# XA1.XA6.MN2.D 0.00176f
C12784 XA6.XA1.XA5.MN2.G D<4> 3.47e-19
C12785 XA5.XA1.XA5.MN2.G XA4.XA6.MN2.D 6.33e-19
C12786 AVDD a_21080_47268# 0.356f
C12787 XA4.XA10.MP0.G VREF 0.0134f
C12788 XDAC1.XC128b<2>.XRES1B.B XDAC1.XC128b<2>.XRES4.B 0.428f
C12789 XB1.XA4.MP0.D m3_n2104_2244# 0.0273f
C12790 a_22448_43748# a_22448_43396# 0.0109f
C12791 XA3.XA1.XA2.MP0.D a_8480_43396# 0.0961f
C12792 XA3.XA1.XA5.MP0.D a_7328_43396# 0.049f
C12793 XA7.XA1.XA2.MP0.D XA7.XA1.XA5.MP0.D 4.34e-19
C12794 SARP XA20.XA1.MN0.D 0.31f
C12795 XA20.XA2a.MN0.D XA6.XA1.XA1.MN0.D 0.0221f
C12796 EN XA7.XA1.XA4.MN1.D 3.17e-19
C12797 XA8.XA1.XA5.MN2.G a_17408_48324# 0.00455f
C12798 XA20.XA10.MN1.D XA20.XA2.MN1.D 0.0138f
C12799 XA3.XA6.MP0.G a_7328_49732# 0.099f
C12800 XA2.XA1.XA5.MN2.G XA0.XA4.MN0.G 6.95e-19
C12801 XA0.XA7.MP0.G XA1.XA4.MN0.G 0.169f
C12802 AVDD XA3.XA1.XA5.MN1.D 0.00889f
C12803 XA7.XA6.MP0.G a_18560_50084# 6.4e-20
C12804 XA7.XA6.MP0.D a_17408_50084# 0.049f
C12805 a_17408_50436# VREF 0.0035f
C12806 XDAC1.XC1.XRES8.B XDAC1.XC1.XRES16.B 0.0904f
C12807 li_9184_7512# li_9184_6900# 0.00271f
C12808 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES1A.B 0.0197f
C12809 XA3.XA3.MN0.G XDAC2.X16ab.XRES16.B 0.00543f
C12810 SARP a_9560_2798# 0.00116f
C12811 XA3.XA1.XA2.MP0.D a_7328_40932# 4.25e-20
C12812 XA1.XA1.XA4.MN0.D a_3440_41988# 0.00176f
C12813 XA6.XA1.XA4.MP0.D a_16040_42340# 0.049f
C12814 a_3440_42340# a_4808_42340# 8.89e-19
C12815 EN a_17408_40228# 0.0658f
C12816 XA20.XA3.MN6.D a_23600_46916# 4.93e-19
C12817 a_9848_48676# a_9848_48324# 0.0109f
C12818 D<7> XA1.XA1.XA5.MN2.D 0.0285f
C12819 XA8.XA7.MP0.G a_19928_45156# 1.95e-19
C12820 XA2.XA1.XA5.MN2.G a_2288_44804# 0.00486f
C12821 XA0.XA7.MP0.G a_3440_44804# 1.95e-19
C12822 AVDD a_21080_41636# 0.404f
C12823 XA5.XA4.MN0.D a_12368_47620# 0.00498f
C12824 VREF a_18560_47620# 7.12e-19
C12825 a_13520_53956# XA6.XA11.MN1.G 0.0225f
C12826 a_12368_53956# XA5.XA12.MP0.G 0.0674f
C12827 AVDD a_5960_53252# 0.364f
C12828 XA0.XA12.MP0.D XA0.XA12.MP0.G 0.142f
C12829 XA20.XA12.MP0.G XA8.XA11.MP0.D 5.54e-19
C12830 a_920_53956# a_920_53604# 0.0109f
C12831 XA1.XA1.XA1.MN0.D a_2288_40932# 8.29e-20
C12832 SARP li_9184_12636# 0.00103f
C12833 VREF a_7328_44100# 0.0251f
C12834 XA2.XA4.MN0.D a_4808_44100# 9.25e-20
C12835 XA20.XA3a.MN0.D a_23600_46212# 8.07e-19
C12836 XA3.XA6.MP0.G XA3.XA1.XA5.MP0.D 0.00121f
C12837 AVDD a_14960_686# 0.37f
C12838 XA0.XA6.MP2.G a_920_42692# 7.76e-20
C12839 XA4.XA1.XA5.MN2.G XA3.XA1.XA4.MN0.D 7.72e-19
C12840 XA5.XA10.MP0.D XA5.XA9.MN1.G 0.00406f
C12841 XA7.XA10.MP0.G XA8.XA10.MP0.G 0.00217f
C12842 a_3440_52900# XA1.XA9.MN1.G 0.00113f
C12843 XA20.XA10.MN1.D a_23600_51844# 0.00466f
C12844 CK_SAMPLE a_n232_51140# 0.0686f
C12845 AVDD D<4> 2.31f
C12846 D<8> a_n232_43748# 0.00363f
C12847 XA1.XA4.MN0.G XA1.XA1.XA4.MP1.D 0.0488f
C12848 XA20.XA3a.MN0.D a_17408_43396# 0.00213f
C12849 CK_SAMPLE a_4808_48676# 4.46e-19
C12850 AVDD a_19928_48324# 0.00166f
C12851 a_8480_51492# a_9848_51492# 8.89e-19
C12852 XA8.XA9.MN1.G XA8.XA6.MP2.D 0.0618f
C12853 a_16040_53604# VREF 0.00351f
C12854 XA20.XA3a.MN0.D a_16040_40932# 0.0658f
C12855 XA7.XA1.XA5.MN1.D a_18560_43748# 0.0494f
C12856 EN XA3.XA1.XA5.MN0.D 0.0063f
C12857 XA2.XA1.XA5.MN1.D XA2.XA1.XA2.MP0.D 0.0102f
C12858 a_21080_50436# a_22448_50436# 8.89e-19
C12859 XA20.XA10.MN1.D a_22448_46212# 2.14e-19
C12860 AVDD a_23600_45156# 0.00159f
C12861 a_12368_51140# VREF 0.00383f
C12862 D<6> a_5960_49732# 0.0109f
C12863 a_7328_50436# XA3.XA6.MP0.G 0.0678f
C12864 a_17408_50788# XA7.XA6.MP0.G 1.34e-19
C12865 XA8.XA1.XA4.MN1.D a_19928_42692# 0.0474f
C12866 XA8.XA1.XA2.MP0.D a_19928_41988# 0.0568f
C12867 XA4.XA1.XA2.MP0.D a_9848_41636# 0.00316f
C12868 XA0.XA1.XA2.MP0.D XA0.XA1.XA1.MN0.S 2.11e-19
C12869 XA3.XA1.XA4.MP1.D XA3.XA1.XA4.MP0.D 0.0488f
C12870 EN XA0.XA1.XA1.MP1.D 6.68e-19
C12871 D<1> XA2.XA3.MN0.G 0.0298f
C12872 XA2.XA1.XA5.MN2.G a_920_45860# 7.1e-20
C12873 XA0.XA7.MP0.G a_2288_45860# 7.1e-20
C12874 VREF a_17408_48676# 0.0191f
C12875 AVDD XA2.XA1.XA4.MP0.D 0.152f
C12876 D<2> XA5.XA3.MN0.G 1.72e-19
C12877 XA3.XA6.MP0.G a_8480_47620# 4.4e-19
C12878 a_2288_49028# a_3440_49028# 0.00133f
C12879 AVDD a_3440_53956# 0.00166f
C12880 XA20.XA12.MP0.G a_22448_54308# 0.0039f
C12881 XA2.XA1.XA1.MP2.D a_5960_41284# 0.0465f
C12882 a_18560_41636# a_18560_41284# 0.0109f
C12883 XA20.XA3a.MN0.D a_22448_47268# 0.00591f
C12884 XA3.XA4.MN0.G XA4.XA3.MN0.G 0.00211f
C12885 XA4.XA4.MN0.G XA3.XA3.MN0.G 0.0104f
C12886 a_22448_47620# a_23600_47620# 0.00133f
C12887 XA6.XA1.XA5.MN2.G a_14888_43396# 0.00504f
C12888 D<1> a_17408_43748# 7.77e-20
C12889 VREF XA6.XA1.XA5.MN2.D 0.341f
C12890 XA3.XA4.MN0.D XA3.XA1.XA5.MN2.D 0.0264f
C12891 XA20.XA3.MN0.D a_23600_45156# 0.029f
C12892 AVDD a_8408_3502# 0.467f
C12893 XA20.XA3.MN6.D SARP 0.0229f
C12894 XA4.XA11.MN1.G XA3.XA9.MN0.D 1.71e-19
C12895 a_8480_53252# a_8480_52900# 0.0109f
C12896 a_19928_53252# XA8.XA10.MP0.D 0.0692f
C12897 AVDD a_22448_51844# 0.568f
C12898 a_17408_40228# a_17408_39876# 0.0109f
C12899 XA1.XA4.MN0.D a_2288_42692# 9.15e-20
C12900 XA7.XA6.MP0.G a_18560_42340# 7.76e-20
C12901 XA20.XA3a.MN0.D XA4.XA1.XA5.MN1.D 2.15e-19
C12902 a_17408_45860# a_18560_45860# 0.00133f
C12903 D<3> a_12368_41284# 7.77e-20
C12904 XA3.XA6.MP0.G a_8480_41988# 7.76e-20
C12905 XA6.XA4.MN0.G a_16040_43748# 6.3e-19
C12906 XA3.XA3.MN0.G a_7328_44804# 0.00498f
C12907 XA6.XA1.XA5.MN2.G a_13520_40932# 0.00838f
C12908 CK_SAMPLE a_3440_49732# 0.0709f
C12909 a_2288_54308# VREF 0.00579f
C12910 XA5.XA9.MN1.G a_12368_51492# 6.57e-19
C12911 AVDD a_5960_49380# 0.356f
C12912 XA0.XA9.MN1.G XA0.XA7.MP0.G 0.0494f
C12913 XA3.XA7.MP0.D a_7328_51844# 0.133f
C12914 XDAC2.XC0.XRES1B.B XDAC2.XC0.XRES4.B 0.428f
C12915 XA20.XA2a.MN0.D a_8480_42692# 0.00563f
C12916 XA1.XA1.XA5.MN2.D a_3440_43396# 1.28e-19
C12917 XA0.XA4.MN0.D a_920_39876# 9.14e-20
C12918 SARN li_14804_13248# 0.00103f
C12919 a_11000_44100# a_12368_44100# 8.89e-19
C12920 XA0.XA6.MP2.G XDAC1.XC64b<1>.XRES8.B 4.06e-21
C12921 AVDD a_21080_46212# 0.356f
C12922 XA5.XA7.MP0.D VREF 0.0234f
C12923 D<6> a_5960_50436# 0.0879f
C12924 XA2.XA6.MN2.D a_4808_50436# 0.00176f
C12925 D<2> a_16040_50788# 0.161f
C12926 XA6.XA6.MN2.D a_14888_50788# 0.0488f
C12927 a_5960_51140# XA2.XA6.MP0.G 6.76e-20
C12928 XA6.XA1.XA5.MN2.G XA5.XA6.MP0.G 0.185f
C12929 li_14804_17952# li_14804_17340# 0.00271f
C12930 XDAC2.XC128a<1>.XRES8.B XDAC2.XC128a<1>.XRES16.B 0.0904f
C12931 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC32a<0>.XRES1B.B 0.00444f
C12932 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES1A.B 0.0197f
C12933 XA20.XA2a.MN0.D a_4808_39876# 1.09e-19
C12934 a_11000_43044# a_12368_43044# 8.89e-19
C12935 XA0.XA6.MP0.G XDAC2.XC1.XRES8.B 0.00687f
C12936 EN a_9848_41988# 1.25e-19
C12937 a_2288_49732# a_2288_49380# 0.0109f
C12938 a_11000_49732# XA4.XA4.MN0.D 0.0658f
C12939 a_16040_49732# VREF 0.029f
C12940 XA3.XA6.MP0.G a_7328_48676# 0.0881f
C12941 XA8.XA1.XA5.MN2.G a_17408_47268# 0.00363f
C12942 AVDD a_14888_43396# 0.00125f
C12943 XA0.XA7.MP0.G a_920_46916# 0.00455f
C12944 XA7.XA6.MP0.G a_17408_49028# 0.0307f
C12945 a_22448_41988# a_23600_41988# 0.00133f
C12946 a_11000_42340# XA4.XA1.XA1.MN0.S 1.34e-19
C12947 VREF a_19928_46564# 7.39e-19
C12948 XA5.XA4.MN0.D a_13520_46564# 4.06e-19
C12949 AVDD a_13520_40932# 0.00125f
C12950 XA20.XA3.MN6.D a_23600_45860# 0.154f
C12951 XA4.XA1.XA5.MN2.G XA4.XA1.XA5.MN1.D 0.0102f
C12952 AVDD a_18560_52548# 0.00166f
C12953 a_19928_53604# a_21080_53604# 0.00133f
C12954 XA6.XA11.MN1.G a_14888_53252# 0.0689f
C12955 XA5.XA12.MP0.G a_13520_53252# 0.0661f
C12956 a_9848_40580# a_11000_40580# 0.00133f
C12957 XA2.XA4.MN0.G a_5960_44452# 5.54e-19
C12958 XA7.XA1.XA5.MN2.G a_18560_41636# 0.0039f
C12959 XA8.XA1.XA5.MN2.G a_17408_41636# 0.0736f
C12960 XA0.XA7.MP0.G XA0.XA1.XA1.MP2.D 0.0736f
C12961 XA2.XA1.XA5.MN2.G XA0.XA1.XA1.MN0.S 3.84e-21
C12962 XA20.XA3a.MN0.D XA20.XA2.MN1.D 0.0184f
C12963 a_4808_52548# XA2.XA7.MP0.D 5.16e-20
C12964 XA6.XA9.MN1.G XA6.XA9.MN0.D 0.034f
C12965 a_16040_52548# a_16040_52196# 0.0109f
C12966 XA8.XA10.MP0.G XA8.XA7.MP0.D 0.0601f
C12967 XA2.XA10.MP0.G a_5960_51844# 0.00224f
C12968 XA1.XA9.MN0.D a_3440_52196# 0.0492f
C12969 XA1.XA9.MN1.G a_4808_52196# 2.84e-19
C12970 CK_SAMPLE a_3440_50436# 0.161f
C12971 AVDD XA5.XA6.MP0.G 5.95f
C12972 XB2.M1.G CK_SAMPLE_BSSW 0.00269f
C12973 XB1.XA3.MN1.D a_8408_1390# 0.0675f
C12974 XB2.XA3.MN0.S XB2.XA3.MN1.D 0.0944f
C12975 XB1.XA3.MN0.S a_9560_1390# 0.0963f
C12976 XB1.M1.G a_11000_334# 0.157f
C12977 XA4.XA6.MP0.G a_11000_40228# 5.5e-19
C12978 XA0.XA6.MP0.G a_920_39876# 0.00207f
C12979 XA20.XA3a.MN0.D XA3.XA1.XA4.MP0.D 1.1e-19
C12980 XA20.XA2a.MN0.D XA7.XA1.XA2.MP0.D 0.227f
C12981 XA5.XA4.MN0.G a_13520_42340# 7.97e-19
C12982 XA6.XA1.XA5.MN2.D a_16040_44100# 0.126f
C12983 SARN XA20.XA3a.MN0.G 0.0883f
C12984 a_16040_51140# a_17408_51140# 8.89e-19
C12985 XA5.XA1.XA5.MN2.G D<4> 0.627f
C12986 AVDD a_19928_47268# 0.00129f
C12987 XA3.XA10.MP0.G VREF 0.0134f
C12988 XB1.XA4.MP0.D m3_7544_2420# 0.106f
C12989 XA20.XA2a.MN0.D XA5.XA1.XA1.MN0.D 0.022f
C12990 EN XA7.XA1.XA4.MP1.D 0.0386f
C12991 XA8.XA1.XA5.MN2.G a_16040_48324# 7.1e-20
C12992 XA7.XA1.XA5.MN2.G a_17408_48324# 7.1e-20
C12993 D<6> a_5960_48676# 0.00918f
C12994 XA0.XA7.MP0.G XA0.XA4.MN0.G 0.158f
C12995 AVDD XA3.XA1.XA5.MP1.D 0.0889f
C12996 D<2> a_16040_49028# 0.00884f
C12997 XA7.XA6.MP0.G a_17408_50084# 0.159f
C12998 a_2288_50084# a_3440_50084# 0.00133f
C12999 a_16040_50436# VREF 0.0035f
C13000 XA20.XA10.MN1.D a_23600_45156# 0.00517f
C13001 XA2.XA3.MN0.G XDAC2.X16ab.XRES16.B 9.19e-20
C13002 D<8> li_14804_23688# 3.5e-20
C13003 XA6.XA1.XA4.MP0.D a_14888_42340# 2.16e-19
C13004 XA6.XA1.XA4.MN0.D a_16040_42340# 2.16e-19
C13005 EN a_16040_40228# 0.0674f
C13006 XA20.XA3a.MN0.G a_23600_46916# 0.154f
C13007 XA20.XA3.MN6.D a_22448_46916# 0.00916f
C13008 a_21080_48676# a_22448_48676# 8.89e-19
C13009 XA8.XA1.XA5.MN2.G a_19928_45156# 1e-19
C13010 XA0.XA7.MP0.G a_2288_44804# 7.1e-20
C13011 XA2.XA1.XA5.MN2.G a_920_44804# 7.1e-20
C13012 AVDD a_19928_41636# 0.00159f
C13013 VREF a_17408_47620# 0.0671f
C13014 a_12368_53956# XA6.XA11.MN1.G 0.0295f
C13015 AVDD a_4808_53252# 0.00154f
C13016 a_14888_41284# a_14888_40932# 0.0109f
C13017 XA1.XA1.XA1.MP1.D a_2288_40932# 0.0465f
C13018 VREF a_5960_44100# 0.0251f
C13019 XA20.XA3a.MN0.D a_22448_46212# 0.00511f
C13020 XA3.XA6.MP0.G XA3.XA1.XA2.MP0.D 0.0106f
C13021 XA2.XA4.MN0.G a_5960_45508# 6.57e-19
C13022 AVDD a_13808_686# 0.00165f
C13023 a_16040_46916# a_17408_46916# 8.89e-19
C13024 a_5960_46916# XA2.XA3.MN0.G 0.0658f
C13025 XA0.XA6.MP2.G a_n232_42692# 6.49e-19
C13026 XA4.XA1.XA5.MN2.G XA3.XA1.XA4.MP0.D 0.00361f
C13027 XA3.XA1.XA5.MN2.G XA3.XA1.XA4.MN0.D 0.00313f
C13028 AVDD XA3.XA6.MN2.D 3.77e-19
C13029 XA6.XA11.MN1.G XA5.XA8.MP0.D 2.37e-19
C13030 a_14888_52900# a_14888_52548# 0.0109f
C13031 XA1.XA10.MP0.G a_3440_52548# 0.13f
C13032 XA20.XA10.MN1.D a_22448_51844# 1.97e-19
C13033 CK_SAMPLE XA8.XA7.MP0.G 0.0785f
C13034 a_9560_3150# XB1.M1.G 0.00116f
C13035 a_8408_3150# XB1.XA4.MP0.D 0.00252f
C13036 a_11000_2798# SAR_IP 0.00271f
C13037 a_14960_3150# XB2.XA1.MP0.D 4.43e-19
C13038 a_18560_45508# a_18560_45156# 0.0109f
C13039 XA3.XA1.XA5.MN2.D a_8480_45156# 0.153f
C13040 a_n232_45156# a_920_45156# 0.00133f
C13041 XA7.XA4.MN0.G a_18560_43044# 0.0409f
C13042 SARN a_12368_n18# 0.00238f
C13043 XA20.XA3a.MN0.D a_16040_43396# 0.00213f
C13044 XA7.XA7.MP0.D a_18560_51140# 0.00388f
C13045 CK_SAMPLE a_3440_48676# 4.46e-19
C13046 AVDD a_18560_48324# 0.00131f
C13047 XA7.XA8.MP0.D a_18560_51492# 0.00224f
C13048 XA8.XA9.MN1.G XA8.XA6.MN2.D 0.126f
C13049 XDAC1.XC64b<1>.XRES8.B XDAC1.XC64b<1>.XRES1A.B 0.0228f
C13050 XDAC1.XC64b<1>.XRES2.B XDAC1.XC64b<1>.XRES16.B 0.457f
C13051 XA20.XA3a.MN0.D a_14888_40932# 0.0739f
C13052 XA20.XA2a.MN0.D a_22448_41988# 0.00423f
C13053 XA7.XA1.XA5.MN1.D a_17408_43748# 2.16e-19
C13054 XA7.XA1.XA5.MP1.D a_18560_43748# 2.16e-19
C13055 a_5960_43748# a_7328_43748# 8.89e-19
C13056 XA0.XA6.MP2.G li_9184_18564# 0.00508f
C13057 a_14888_44100# XA6.XA1.XA2.MP0.D 2.92e-19
C13058 EN XA3.XA1.XA5.MP0.D 0.0446f
C13059 D<2> a_16040_50084# 0.0155f
C13060 XA4.XA1.XA5.MN2.G a_7328_49380# 0.00363f
C13061 AVDD a_22448_45156# 0.405f
C13062 a_11000_51140# VREF 0.00383f
C13063 D<6> a_4808_49732# 7.01e-19
C13064 XDAC1.XC32a<0>.XRES2.B XDAC1.XC64a<0>.XRES2.B 1.67e-19
C13065 XA0.XA4.MN0.D XDAC1.XC1.XRES8.B 0.00687f
C13066 a_7328_42692# a_8480_42692# 0.00133f
C13067 EN XA0.XA1.XA1.MN0.D 0.0229f
C13068 D<1> XA1.XA3.MN0.G 0.0298f
C13069 XA0.XA7.MP0.G a_920_45860# 0.00363f
C13070 XA4.XA4.MN0.D a_11000_48676# 0.154f
C13071 VREF a_16040_48676# 0.0191f
C13072 AVDD XA2.XA1.XA4.MN0.D 0.00889f
C13073 XA3.XA6.MP0.G a_7328_47620# 6.35e-19
C13074 XA7.XA6.MP0.G a_18560_47972# 6.28e-19
C13075 a_14888_49380# a_14888_49028# 0.0109f
C13076 XA8.XA1.XA5.MN2.G a_17408_46212# 0.00363f
C13077 AVDD a_2288_53956# 0.464f
C13078 XA20.XA12.MP0.D a_22448_54308# 0.0271f
C13079 XA20.XA12.MP0.G a_21080_54308# 0.00424f
C13080 a_22448_55012# CK_SAMPLE 2.89e-19
C13081 a_5960_54308# a_7328_54308# 8.89e-19
C13082 SARP XDAC1.X16ab.XRES1A.B 3.59f
C13083 XA2.XA1.XA1.MN0.S a_5960_41284# 0.0964f
C13084 XA3.XA4.MN0.G XA3.XA3.MN0.G 0.639f
C13085 a_9848_47620# a_9848_47268# 0.0109f
C13086 D<6> XA2.XA1.XA5.MP0.D 7.42e-19
C13087 XA5.XA1.XA5.MN2.G a_14888_43396# 7.1e-20
C13088 XA6.XA1.XA5.MN2.G a_13520_43396# 2.66e-19
C13089 XA1.XA6.MP0.G a_3440_44100# 7.76e-20
C13090 VREF XA5.XA1.XA5.MN2.D 0.341f
C13091 XA20.XA3.MN0.D a_22448_45156# 2.46e-19
C13092 AVDD a_9560_3854# 0.00166f
C13093 XA5.XA6.MP0.G a_13520_44452# 7.76e-20
C13094 XA20.XA3a.MN0.G SARP 2.28e-19
C13095 XA20.XA3.MN6.D a_23600_44804# 0.068f
C13096 XA4.XA11.MN1.G XA3.XA9.MN1.G 0.0169f
C13097 XA1.XA10.MP0.D XA2.XA10.MP0.D 0.00217f
C13098 AVDD a_21080_51844# 0.385f
C13099 a_19928_53956# XA8.XA9.MN1.G 7.37e-20
C13100 a_3440_39876# a_4808_39876# 8.89e-19
C13101 XA7.XA6.MP0.G a_17408_42340# 5.5e-19
C13102 XA20.XA3a.MN0.D XA3.XA1.XA5.MN1.D 2.15e-19
C13103 a_4808_45860# a_4808_45508# 0.0109f
C13104 XA3.XA6.MP0.G a_7328_41988# 5.5e-19
C13105 XA6.XA4.MN0.G a_14888_43748# 0.0157f
C13106 XA5.XA1.XA5.MN2.G a_13520_40932# 0.00631f
C13107 XA6.XA1.XA5.MN2.G a_12368_40932# 0.0245f
C13108 CK_SAMPLE a_2288_49732# 0.00347f
C13109 a_920_54308# VREF 0.00579f
C13110 AVDD a_4808_49380# 0.00159f
C13111 a_16040_52548# XA7.XA1.XA5.MN2.G 1.75e-19
C13112 a_17408_52196# a_17408_51844# 0.0109f
C13113 a_n232_44804# XA0.XA1.XA2.MP0.D 2.6e-20
C13114 XA20.XA2a.MN0.D a_7328_42692# 0.00457f
C13115 XA1.XA1.XA5.MN2.D a_2288_43396# 4.58e-19
C13116 D<7> XDAC1.XC64b<1>.XRES4.B 0.00405f
C13117 XA0.XA4.MN0.D a_n232_39876# 9.25e-20
C13118 a_23600_44452# a_23600_44100# 0.0109f
C13119 AVDD a_19928_46212# 0.00154f
C13120 a_920_50788# a_2288_50788# 8.89e-19
C13121 XA4.XA7.MP0.D VREF 0.0234f
C13122 D<6> a_4808_50436# 5.7e-19
C13123 XA5.XA1.XA5.MN2.G XA5.XA6.MP0.G 0.0738f
C13124 XA20.XA2a.MN0.D a_3440_39876# 1.09e-19
C13125 a_23600_43396# a_23600_43044# 0.0109f
C13126 EN a_8480_41988# 1.25e-19
C13127 a_9848_49732# XA4.XA4.MN0.D 0.0675f
C13128 a_19928_49732# a_21080_49732# 0.00133f
C13129 D<4> XA20.XA3a.MN0.D 0.0799f
C13130 D<6> a_5960_47620# 0.0147f
C13131 XA7.XA1.XA5.MN2.G a_17408_47268# 7.1e-20
C13132 XA8.XA1.XA5.MN2.G a_16040_47268# 7.1e-20
C13133 AVDD a_13520_43396# 0.00125f
C13134 a_9848_41988# a_9848_41636# 0.0109f
C13135 VREF a_18560_46564# 7.39e-19
C13136 XA5.XA4.MN0.D a_12368_46564# 1.28e-19
C13137 a_3440_47972# a_4808_47972# 8.89e-19
C13138 AVDD a_12368_40932# 0.358f
C13139 XA5.XA6.MP0.G a_13520_45508# 7.76e-20
C13140 XA20.XA3.MN6.D a_22448_45860# 0.164f
C13141 XA5.XA4.MN0.G a_13520_47972# 0.153f
C13142 a_22448_48324# a_22448_47972# 0.0109f
C13143 XA4.XA1.XA5.MN2.G XA3.XA1.XA5.MN1.D 6.68e-19
C13144 XA0.XA12.MP0.G XA0.XA10.MP0.D 0.0632f
C13145 XA0.XA12.MP0.D XA1.XA10.MP0.D 0.0909f
C13146 AVDD a_17408_52548# 0.405f
C13147 a_920_53604# a_920_53252# 0.0109f
C13148 XA5.XA12.MP0.G a_12368_53252# 0.00276f
C13149 XA6.XA11.MN1.G a_13520_53252# 0.0238f
C13150 a_22448_40932# a_22448_40580# 0.0109f
C13151 a_11000_46564# a_11000_46212# 0.0109f
C13152 a_23600_46564# XA20.XA2a.MN0.D 0.00238f
C13153 XA2.XA3.MN0.G a_5960_45860# 0.155f
C13154 XA2.XA4.MN0.G a_4808_44452# 0.00907f
C13155 D<6> a_5960_41988# 7.76e-20
C13156 XA7.XA1.XA5.MN2.G a_17408_41636# 4.13e-19
C13157 XA0.XA11.MN1.G a_13808_1742# 0.00212f
C13158 XA0.XA7.MP0.G XA0.XA1.XA1.MN0.S 0.327f
C13159 XA4.XA6.MP0.G XA4.XA1.XA4.MP1.D 0.00121f
C13160 VREF XA5.XA1.XA5.MP0.D 0.00202f
C13161 D<2> a_16040_42340# 7.76e-20
C13162 XA2.XA10.MP0.G a_4808_51844# 5.59e-19
C13163 XA1.XA9.MN1.G a_3440_52196# 0.0878f
C13164 CK_SAMPLE a_2288_50436# 0.00312f
C13165 AVDD XA4.XA6.MP0.D 0.144f
C13166 XB2.M1.G a_14960_686# 8.55e-20
C13167 SAR_IN a_12368_n18# 0.0347f
C13168 XB1.XA4.MP0.D a_8408_334# 0.00258f
C13169 XB1.XA3.MN0.S a_8408_1390# 1.28e-19
C13170 a_12368_1742# a_12368_1390# 0.0109f
C13171 SARN li_14804_23688# 0.00103f
C13172 XA2.XA4.MN0.D XA2.XA1.XA1.MN0.D 0.00301f
C13173 XA4.XA6.MP0.G a_9848_40228# 7.76e-20
C13174 XA0.XA6.MP0.G a_n232_39876# 7.76e-20
C13175 XA20.XA3a.MN0.D XA2.XA1.XA4.MP0.D 1.1e-19
C13176 a_17408_44804# a_18560_44804# 0.00133f
C13177 a_4808_44804# a_4808_44452# 0.0109f
C13178 XA5.XA4.MN0.G a_12368_42340# 1.28e-19
C13179 XA7.XA3.MN0.G a_18560_43396# 6.8e-20
C13180 XA6.XA1.XA5.MN2.D a_14888_44100# 0.0877f
C13181 a_2288_51140# XA1.XA6.MP2.D 0.00176f
C13182 XA4.XA1.XA5.MN2.G D<4> 0.00595f
C13183 AVDD a_18560_47268# 0.00125f
C13184 a_17408_51492# D<1> 2.41e-19
C13185 XA2.XA10.MP0.G VREF 0.0134f
C13186 XDAC2.X16ab.XRES2.B XDAC2.XC128b<2>.XRES2.B 1.67e-19
C13187 li_14804_23076# li_14804_22656# 0.00411f
C13188 XB1.XA4.MP0.D m3_7472_2420# 0.0634f
C13189 a_21080_43748# a_21080_43396# 0.0109f
C13190 XA20.XA2a.MN0.D XA5.XA1.XA1.MP1.D 0.00946f
C13191 EN XA6.XA1.XA4.MP1.D 0.0386f
C13192 XA7.XA1.XA5.MN2.G a_16040_48324# 0.00455f
C13193 D<6> a_4808_48676# 3.48e-19
C13194 XA2.XA6.MP0.D a_5960_49732# 0.00176f
C13195 D<2> a_14888_49028# 5.7e-19
C13196 AVDD XA2.XA1.XA5.MP1.D 0.0889f
C13197 XA20.XA10.MN1.D a_22448_45156# 2.14e-19
C13198 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES1A.B 0.00438f
C13199 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES16.B 0.0483f
C13200 XDAC2.XC1.XRES8.B XDAC2.XC1.XRES2.B 0.44f
C13201 XA3.XA3.MN0.G li_14804_24300# 0.00504f
C13202 XA1.XA1.XA4.MP0.D a_2288_41988# 0.00176f
C13203 XA6.XA1.XA4.MN0.D a_14888_42340# 0.0474f
C13204 a_2288_42340# a_3440_42340# 0.00133f
C13205 XA20.XA3a.MN0.G a_22448_46916# 0.183f
C13206 XA3.XA6.MP0.G a_8480_46564# 7.76e-20
C13207 a_8480_48676# a_8480_48324# 0.0109f
C13208 XA8.XA1.XA5.MN2.G a_18560_45156# 1.95e-19
C13209 XA0.XA7.MP0.G a_920_44804# 0.00486f
C13210 AVDD a_18560_41636# 0.00125f
C13211 VREF a_16040_47620# 0.0671f
C13212 XA4.XA4.MN0.D a_11000_47620# 0.00498f
C13213 AVDD a_3440_53252# 0.00144f
C13214 a_13520_53956# XA5.XA11.MN1.G 0.00258f
C13215 a_n232_53956# a_n232_53604# 0.0109f
C13216 XA5.XA1.XA1.MN0.S a_13520_40580# 0.00155f
C13217 XA0.XA1.XA1.MN0.S a_920_40228# 0.0313f
C13218 SARP li_9184_13248# 0.00103f
C13219 XA1.XA4.MN0.D a_3440_44100# 9.24e-20
C13220 XA2.XA4.MN0.G a_4808_45508# 0.0104f
C13221 a_4808_46916# XA2.XA3.MN0.G 0.0682f
C13222 XA3.XA1.XA5.MN2.G XA3.XA1.XA4.MP0.D 6.33e-19
C13223 AVDD XA3.XA6.MP2.D 0.172f
C13224 XA1.XA10.MP0.G a_2288_52548# 0.0684f
C13225 XA6.XA10.MP0.G XA7.XA10.MP0.G 0.00217f
C13226 CK_SAMPLE XA8.XA1.XA5.MN2.G 0.0595f
C13227 a_8408_3150# XB1.M1.G 2.71e-20
C13228 XB1.XA2.MN0.G XB1.XA4.MP0.D 0.0112f
C13229 a_13808_2798# a_14960_2798# 0.00133f
C13230 a_13808_3150# XB2.XA1.MP0.D 0.00203f
C13231 XA3.XA1.XA5.MN2.D a_7328_45156# 0.155f
C13232 XA7.XA4.MN0.G a_17408_43044# 0.0222f
C13233 XA0.XA4.MN0.G XA0.XA1.XA4.MP1.D 0.0488f
C13234 XA8.XA7.MP0.G a_21080_39876# 0.00141f
C13235 D<1> a_18560_40580# 5.26e-19
C13236 D<5> a_8480_40228# 2.88e-19
C13237 SARN a_11000_n18# 1.62e-20
C13238 XA20.XA3a.MN0.D a_14888_43396# 0.0736f
C13239 a_17408_51844# XA8.XA1.XA5.MN2.G 8.87e-19
C13240 XA7.XA7.MP0.D a_17408_51140# 0.00224f
C13241 CK_SAMPLE a_2288_48676# 6.2e-20
C13242 AVDD a_17408_48324# 0.359f
C13243 XA8.XA9.MN1.G D<0> 0.0378f
C13244 a_7328_51492# a_8480_51492# 0.00133f
C13245 XA7.XA8.MP0.D a_17408_51492# 0.00224f
C13246 XA3.XA9.MN1.G a_8480_50788# 0.015f
C13247 a_11000_52196# D<4> 7.56e-20
C13248 XA20.XA3a.MN0.D a_13520_40932# 0.0723f
C13249 XA5.XA1.XA5.MN2.D a_12368_42692# 7.44e-20
C13250 XA20.XA2a.MN0.D a_21080_41988# 0.0044f
C13251 XA7.XA1.XA5.MP1.D a_17408_43748# 0.049f
C13252 XA2.XA3.MN0.G XA2.XA1.XA1.MN0.S 0.0101f
C13253 XA1.XA1.XA5.MN1.D XA1.XA1.XA5.MN0.D 0.0488f
C13254 EN XA3.XA1.XA2.MP0.D 0.03f
C13255 D<2> a_14888_50084# 5.7e-19
C13256 a_19928_50436# a_21080_50436# 0.00133f
C13257 XA3.XA1.XA5.MN2.G a_7328_49380# 7.1e-20
C13258 XA4.XA1.XA5.MN2.G a_5960_49380# 7.1e-20
C13259 AVDD a_21080_45156# 0.356f
C13260 a_5960_50436# XA2.XA6.MP0.D 0.00176f
C13261 XA7.XA1.XA4.MN1.D a_18560_42692# 0.0474f
C13262 XA2.XA1.XA4.MP1.D XA2.XA1.XA4.MP0.D 0.0488f
C13263 AVDD XA1.XA1.XA4.MN0.D 0.00889f
C13264 D<1> D<8> 0.0362f
C13265 VREF a_14888_48676# 1.3e-19
C13266 XA4.XA4.MN0.D a_9848_48676# 0.158f
C13267 XA5.XA6.MP0.G XA20.XA3a.MN0.D 0.0759f
C13268 D<2> XA3.XA3.MN0.G 0.0319f
C13269 D<3> XA6.XA3.MN0.G 1.72e-19
C13270 D<0> a_21080_46916# 0.0185f
C13271 XA7.XA6.MP0.G a_17408_47972# 8.92e-19
C13272 a_920_49028# a_2288_49028# 8.89e-19
C13273 XA7.XA1.XA5.MN2.G a_17408_46212# 7.1e-20
C13274 XA8.XA1.XA5.MN2.G a_16040_46212# 7.1e-20
C13275 AVDD a_920_53956# 0.461f
C13276 XA20.XA12.MP0.G a_19928_54308# 2.54e-19
C13277 XA6.XA1.XA1.MN0.S XA7.XA1.XA1.MN0.S 0.00217f
C13278 XA2.XA1.XA1.MN0.S a_4808_41284# 0.0658f
C13279 a_17408_41636# a_17408_41284# 0.0109f
C13280 XA8.XA4.MN0.G a_21080_46916# 0.0678f
C13281 a_21080_47620# a_22448_47620# 8.89e-19
C13282 D<6> XA2.XA1.XA5.MN0.D 0.00188f
C13283 XA5.XA1.XA5.MN2.G a_13520_43396# 0.00518f
C13284 XA6.XA1.XA5.MN2.G a_12368_43396# 0.00442f
C13285 XA1.XA6.MP0.G a_2288_44100# 5.5e-19
C13286 VREF XA4.XA1.XA5.MN2.D 0.341f
C13287 XA2.XA4.MN0.D XA2.XA1.XA5.MN2.D 0.0265f
C13288 AVDD a_8408_3854# 0.448f
C13289 XA5.XA6.MP0.G a_12368_44452# 5.5e-19
C13290 XA20.XA3a.MN0.G a_23600_44804# 0.00276f
C13291 XA20.XA3.MN6.D a_22448_44804# 0.174f
C13292 a_7328_53252# a_7328_52900# 0.0109f
C13293 a_18560_53252# XA7.XA10.MP0.D 0.0676f
C13294 XA7.XA11.MP0.D a_17408_52900# 0.00176f
C13295 AVDD a_19928_51844# 0.00166f
C13296 XA3.XA11.MN1.G XA3.XA9.MN0.D 1.35e-19
C13297 a_16040_40228# a_16040_39876# 0.0109f
C13298 SARN a_13808_3150# 0.00116f
C13299 XA20.XA3a.MN0.D XA3.XA1.XA5.MP1.D 2.15e-19
C13300 a_16040_45860# a_17408_45860# 8.89e-19
C13301 XA2.XA3.MN0.G a_5960_44804# 0.00498f
C13302 XA5.XA1.XA5.MN2.G a_12368_40932# 0.0013f
C13303 CK_SAMPLE a_920_49732# 0.00347f
C13304 AVDD a_3440_49380# 0.00159f
C13305 XA2.XA7.MP0.D a_5960_51844# 0.133f
C13306 XDAC1.XC0.XRES1B.B XDAC1.XC0.XRES4.B 0.428f
C13307 XA20.XA2a.MN0.D a_5960_42692# 0.00457f
C13308 a_9848_45156# XA4.XA1.XA2.MP0.D 1.56e-20
C13309 XA0.XA6.MP2.G li_9184_29004# 3.5e-20
C13310 SARN XDAC2.XC32a<0>.XRES16.B 55.3f
C13311 a_9848_44100# a_11000_44100# 0.00133f
C13312 a_21080_44452# EN 0.00173f
C13313 XA20.XA3a.MN0.D a_19928_41636# 0.00547f
C13314 AVDD a_18560_46212# 0.00125f
C13315 XA8.XA9.MN1.G a_21080_49380# 2.54e-19
C13316 XA3.XA7.MP0.D VREF 0.0234f
C13317 XDAC1.XC128a<1>.XRES8.B XDAC1.XC128a<1>.XRES16.B 0.0904f
C13318 li_9184_17952# li_9184_17340# 0.00271f
C13319 XDAC1.XC128a<1>.XRES1B.B XDAC1.XC32a<0>.XRES1B.B 0.00444f
C13320 XDAC1.XC128a<1>.XRES4.B XDAC1.XC128a<1>.XRES1A.B 0.0197f
C13321 XA1.XA1.XA2.MP0.D XA1.XA1.XA4.MN0.D 0.056f
C13322 XA5.XA1.XA2.MP0.D a_13520_42692# 0.0946f
C13323 a_9848_43044# a_11000_43044# 0.00133f
C13324 XA0.XA6.MP0.G li_14804_8124# 0.00506f
C13325 EN a_7328_41988# 0.0723f
C13326 D<6> a_4808_47620# 5.21e-19
C13327 XA7.XA1.XA5.MN2.G a_16040_47268# 0.00363f
C13328 D<2> a_16040_47972# 0.0147f
C13329 AVDD a_12368_43396# 0.361f
C13330 a_920_49732# a_920_49380# 0.0109f
C13331 a_21080_41988# a_22448_41988# 8.89e-19
C13332 SARP a_11000_n18# 0.00258f
C13333 AVDD a_11000_40932# 0.358f
C13334 VREF a_17408_46564# 0.0175f
C13335 XA5.XA6.MP0.G a_12368_45508# 5.5e-19
C13336 XA0.XA6.MP2.G a_920_44100# 7.76e-20
C13337 XA20.XA3a.MN0.G a_22448_45860# 0.0277f
C13338 XA5.XA4.MN0.G a_12368_47972# 0.155f
C13339 XA3.XA1.XA5.MN2.G XA3.XA1.XA5.MN1.D 0.0102f
C13340 XA4.XA1.XA5.MN2.G XA3.XA1.XA5.MP1.D 0.00329f
C13341 D<4> a_11000_44452# 1.47e-19
C13342 XA0.XA12.MP0.D XA0.XA10.MP0.D 0.00744f
C13343 XA5.XA11.MN1.G a_14888_53252# 2.81e-19
C13344 a_18560_53604# a_19928_53604# 8.89e-19
C13345 XA6.XA11.MN1.G a_12368_53252# 3.16e-19
C13346 AVDD a_16040_52548# 0.405f
C13347 a_8480_40580# a_9848_40580# 8.89e-19
C13348 a_22448_46564# XA20.XA2a.MN0.D 0.00224f
C13349 XA2.XA3.MN0.G a_4808_45860# 0.162f
C13350 XA2.XA4.MN0.G a_3440_44452# 2.2e-19
C13351 XA1.XA4.MN0.G a_4808_44452# 2.2e-19
C13352 D<6> a_4808_41988# 6.49e-19
C13353 XA7.XA1.XA5.MN2.G a_16040_41636# 0.0756f
C13354 XA0.XA11.MN1.G a_12368_1742# 0.156f
C13355 XA4.XA6.MP0.G XA4.XA1.XA4.MN1.D 7.41e-19
C13356 D<2> a_14888_42340# 6.49e-19
C13357 XA20.XA3a.MN0.D a_22448_45156# 0.00524f
C13358 a_3440_52548# XA1.XA7.MP0.D 5.16e-20
C13359 XA7.XA10.MP0.G XA7.XA7.MP0.D 0.0601f
C13360 AVDD XA4.XA6.MN0.D 3.13e-19
C13361 a_14888_52548# a_14888_52196# 0.0109f
C13362 XA1.XA9.MN1.G a_2288_52196# 0.0665f
C13363 CK_SAMPLE a_920_50436# 0.00312f
C13364 XB1.XA4.MP0.D CK_SAMPLE_BSSW 0.00524f
C13365 XB1.M1.G a_8408_334# 3.51e-20
C13366 XB1.XA0.MP0.D a_9560_1038# 0.158f
C13367 XA20.XA3a.MN0.D XA2.XA1.XA4.MN0.D 1.1e-19
C13368 a_21080_45508# EN 1.42e-19
C13369 XA4.XA1.XA5.MN2.G XA3.XA6.MN2.D 6.33e-19
C13370 XA3.XA9.MN1.G a_8480_50084# 0.00969f
C13371 XA8.XA7.MP0.D a_19928_50436# 1.37e-19
C13372 a_2288_51140# D<7> 0.0688f
C13373 a_14888_51140# a_16040_51140# 0.00133f
C13374 XA3.XA1.XA5.MN2.G D<4> 4.48e-21
C13375 AVDD a_17408_47268# 0.356f
C13376 XA1.XA10.MP0.G VREF 0.0134f
C13377 XB1.XA4.MP0.D m3_n1960_3300# 0.0137f
C13378 XA2.XA1.XA5.MP0.D a_5960_43396# 0.049f
C13379 XA20.XA2a.MN0.D XA4.XA1.XA1.MP1.D 0.00946f
C13380 D<8> a_n232_40580# 0.00369f
C13381 EN XA6.XA1.XA4.MN1.D 3.17e-19
C13382 AVDD XA2.XA1.XA5.MN1.D 0.00889f
C13383 XA6.XA6.MP0.D a_16040_50084# 0.049f
C13384 a_920_50084# a_2288_50084# 8.89e-19
C13385 D<8> XDAC2.X16ab.XRES16.B 3.84e-19
C13386 D<0> a_21080_45860# 0.0777f
C13387 a_19928_48676# a_21080_48676# 0.00133f
C13388 XA6.XA6.MP0.G XA6.XA3.MN0.G 0.0501f
C13389 XA3.XA6.MP0.G a_7328_46564# 5.5e-19
C13390 D<4> a_11000_45508# 0.00436f
C13391 XA8.XA1.XA5.MN2.G a_17408_45156# 0.00486f
C13392 XA7.XA1.XA5.MN2.G a_18560_45156# 1e-19
C13393 XA0.XA7.MP0.G a_n232_44804# 1.86e-19
C13394 AVDD a_17408_41636# 0.404f
C13395 XA7.XA6.MP0.G XA3.XA3.MN0.G 0.0371f
C13396 XA4.XA4.MN0.D a_9848_47620# 0.0396f
C13397 VREF a_14888_47620# 7.12e-19
C13398 a_n232_54308# XA0.XA11.MN1.G 2.9e-19
C13399 AVDD a_2288_53252# 0.361f
C13400 a_11000_53956# XA4.XA12.MP0.G 0.0658f
C13401 a_12368_53956# XA5.XA11.MN1.G 0.00198f
C13402 a_13520_41284# a_13520_40932# 0.0109f
C13403 XA0.XA1.XA1.MP1.D a_920_40932# 0.0465f
C13404 XA5.XA1.XA1.MN0.S a_12368_40580# 0.0318f
C13405 XA0.XA1.XA1.MN0.S a_n232_40228# 0.0215f
C13406 XA7.XA6.MP0.G a_18560_43748# 7.76e-20
C13407 D<5> XA3.XA1.XA4.MN1.D 0.00188f
C13408 XA1.XA4.MN0.D a_2288_44100# 9.15e-20
C13409 XA1.XA4.MN0.G a_4808_45508# 2.84e-19
C13410 XA2.XA4.MN0.G a_3440_45508# 2.84e-19
C13411 XA8.XA4.MN0.G a_21080_45860# 2.12e-19
C13412 a_14888_46916# a_16040_46916# 0.00133f
C13413 XA3.XA1.XA5.MN2.G XA2.XA1.XA4.MP0.D 0.00361f
C13414 D<1> a_18560_43044# 6.49e-19
C13415 AVDD D<5> 2.23f
C13416 a_19928_53252# XA8.XA9.MN1.G 5.25e-19
C13417 XA5.XA11.MN1.G XA5.XA8.MP0.D 6.42e-19
C13418 XA4.XA10.MP0.D XA4.XA9.MN1.G 0.00406f
C13419 a_13520_52900# a_13520_52548# 0.0109f
C13420 CK_SAMPLE XA7.XA1.XA5.MN2.G 0.0595f
C13421 XB1.XA2.MN0.G XB1.M1.G 0.00145f
C13422 a_9560_2798# XB1.XA1.MN0.D 0.0958f
C13423 XB2.XA2.MN0.G XB2.XA1.MP0.D 0.00383f
C13424 a_17408_45508# a_17408_45156# 0.0109f
C13425 XA0.XA4.MN0.G XA0.XA1.XA4.MN1.D 0.0642f
C13426 XA1.XA6.MP0.G XA1.XA1.XA1.MN0.D 0.00112f
C13427 D<1> a_17408_40580# 4.18e-20
C13428 D<5> a_7328_40228# 3.45e-20
C13429 XA5.XA6.MP0.G a_13520_41284# 3.97e-20
C13430 XA20.XA3a.MN0.D a_13520_43396# 0.0723f
C13431 XA0.XA7.MP0.D XA0.XA6.MP2.G 2.65e-19
C13432 CK_SAMPLE a_920_48676# 6.2e-20
C13433 AVDD a_16040_48324# 0.359f
C13434 XA3.XA9.MN1.G a_7328_50788# 0.00281f
C13435 SARN D<1> 0.0307f
C13436 a_12368_53604# VREF 0.00396f
C13437 XDAC2.XC64b<1>.XRES8.B XDAC2.XC64b<1>.XRES16.B 0.0904f
C13438 XDAC2.XC64b<1>.XRES1B.B XDAC2.X16ab.XRES1B.B 0.00444f
C13439 XDAC2.XC64b<1>.XRES4.B XDAC2.XC64b<1>.XRES1A.B 0.0197f
C13440 li_14804_28392# li_14804_27780# 0.00271f
C13441 XA20.XA3a.MN0.D a_12368_40932# 0.0674f
C13442 XA20.XA2a.MN0.D a_19928_41988# 0.0851f
C13443 a_4808_43748# a_5960_43748# 0.00133f
C13444 XA0.XA6.MP2.G XDAC1.XC128a<1>.XRES4.B 0.00406f
C13445 XA1.XA3.MN0.G XA2.XA1.XA1.MN0.S 1.07e-19
C13446 EN XA2.XA1.XA5.MP0.D 0.0446f
C13447 XA3.XA1.XA5.MN2.G a_5960_49380# 0.00363f
C13448 AVDD a_19928_45156# 0.00159f
C13449 XA8.XA7.MP0.G XA8.XA4.MN0.D 0.0939f
C13450 li_9184_12636# li_9184_12216# 0.00411f
C13451 a_5960_42692# a_7328_42692# 8.89e-19
C13452 XA7.XA1.XA4.MP1.D a_18560_42692# 2.16e-19
C13453 XA7.XA1.XA4.MN1.D a_17408_42692# 2.16e-19
C13454 EN a_22448_41284# 5.7e-20
C13455 XA0.XA4.MN0.D li_9184_8124# 0.00506f
C13456 AVDD XA1.XA1.XA4.MP0.D 0.152f
C13457 VREF a_13520_48676# 1.3e-19
C13458 D<2> XA2.XA3.MN0.G 0.0309f
C13459 D<3> XA5.XA3.MN0.G 0.572f
C13460 D<0> a_19928_46916# 0.00249f
C13461 a_13520_49380# a_13520_49028# 0.0109f
C13462 D<6> a_5960_46564# 0.0695f
C13463 XA7.XA1.XA5.MN2.G a_16040_46212# 0.00363f
C13464 AVDD a_n232_53956# 0.00164f
C13465 a_22448_55364# CK_SAMPLE 1.64e-19
C13466 a_4808_54308# a_5960_54308# 0.00133f
C13467 SARP li_9184_23688# 0.00103f
C13468 XA6.XA1.XA1.MN0.S XA6.XA1.XA1.MP2.D 0.0708f
C13469 XA8.XA4.MN0.G a_19928_46916# 0.0869f
C13470 XA2.XA4.MN0.G XA2.XA3.MN0.G 0.622f
C13471 a_8480_47620# a_8480_47268# 0.0109f
C13472 D<6> XA2.XA1.XA2.MP0.D 0.0131f
C13473 VREF XA3.XA1.XA5.MN2.D 0.341f
C13474 AVDD a_23600_39876# 0.00148f
C13475 XA20.XA3a.MN0.G a_22448_44804# 0.0724f
C13476 XA0.XA10.MP0.D XA1.XA10.MP0.D 0.00217f
C13477 a_17408_53252# XA7.XA10.MP0.D 0.0677f
C13478 XA8.XA11.MN1.G a_19928_52548# 2.85e-19
C13479 AVDD a_18560_51844# 0.00166f
C13480 XA3.XA11.MN1.G XA3.XA9.MN1.G 0.00349f
C13481 a_2288_39876# a_3440_39876# 0.00133f
C13482 XA0.XA4.MN0.D a_920_42692# 9.14e-20
C13483 SARN XB2.XA2.MN0.G 0.00236f
C13484 XA20.XA2a.MN0.D XA7.XA1.XA5.MN2.D 8.92e-20
C13485 a_3440_45860# a_3440_45508# 0.0109f
C13486 XA5.XA4.MN0.G a_13520_43748# 0.0157f
C13487 XA2.XA3.MN0.G a_4808_44804# 0.043f
C13488 XA20.XA3a.MN0.D XA2.XA1.XA5.MP1.D 2.15e-19
C13489 XA5.XA1.XA5.MN2.G a_11000_40932# 0.0256f
C13490 CK_SAMPLE a_n232_49732# 0.0693f
C13491 AVDD a_2288_49380# 0.356f
C13492 a_4808_52196# XA2.XA8.MP0.D 2.11e-19
C13493 XA20.XA11.MP0.D VREF 2.19e-19
C13494 XA4.XA9.MN1.G a_11000_51492# 6.57e-19
C13495 a_16040_52196# a_16040_51844# 0.0109f
C13496 XA2.XA7.MP0.D a_4808_51844# 0.159f
C13497 XA7.XA7.MP0.D XA8.XA7.MP0.D 0.00435f
C13498 XA20.XA2.MN1.D a_23600_43748# 0.0137f
C13499 XA20.XA2a.MN0.D a_4808_42692# 0.00563f
C13500 XA0.XA1.XA5.MN2.D a_920_43396# 4.58e-19
C13501 XA7.XA1.XA5.MN2.D XA7.XA1.XA2.MP0.D 4.72e-19
C13502 XA8.XA4.MN0.G XA8.XA1.XA1.MN0.S 5.22e-20
C13503 D<7> li_9184_29616# 0.00504f
C13504 a_22448_44452# a_22448_44100# 0.0109f
C13505 a_19928_44452# EN 0.00154f
C13506 XA20.XA3a.MN0.D a_18560_41636# 0.00547f
C13507 AVDD a_17408_46212# 0.356f
C13508 XA6.XA1.XA5.MN2.G XA4.XA6.MP0.G 3.47e-19
C13509 a_n232_50788# a_920_50788# 0.00133f
C13510 XA8.XA9.MN1.G a_19928_49380# 4.23e-20
C13511 XA2.XA7.MP0.D VREF 0.0234f
C13512 XA1.XA6.MN2.D a_3440_50436# 0.00176f
C13513 XA5.XA6.MN2.D a_13520_50788# 0.0488f
C13514 XA5.XA1.XA2.MP0.D a_12368_42692# 7.68e-20
C13515 XA1.XA1.XA2.MP0.D XA1.XA1.XA4.MP0.D 4.34e-19
C13516 a_22448_43396# a_22448_43044# 0.0109f
C13517 EN a_5960_41988# 0.0739f
C13518 D<2> a_14888_47972# 5.43e-19
C13519 AVDD a_11000_43396# 0.361f
C13520 a_18560_49732# a_19928_49732# 8.89e-19
C13521 a_12368_49732# VREF 0.029f
C13522 a_8480_49732# XA3.XA4.MN0.D 0.0659f
C13523 a_8480_41988# a_8480_41636# 0.0109f
C13524 AVDD a_9848_40932# 0.00125f
C13525 VREF a_16040_46564# 0.0175f
C13526 XA4.XA4.MN0.D a_11000_46564# 1.28e-19
C13527 XA0.XA6.MP2.G a_n232_44100# 6.49e-19
C13528 a_2288_47972# a_3440_47972# 0.00133f
C13529 a_21080_48324# a_21080_47972# 0.0109f
C13530 D<0> a_21080_44804# 1.95e-19
C13531 XA1.XA6.MP0.G XA1.XA1.XA5.MN2.D 0.0267f
C13532 XA3.XA1.XA5.MN2.G XA3.XA1.XA5.MP1.D 5.21e-20
C13533 D<4> a_9848_44452# 5.24e-19
C13534 D<1> SARP 0.0443f
C13535 XA5.XA11.MN1.G a_13520_53252# 0.0758f
C13536 a_7328_53604# XA3.XA11.MP0.D 0.00176f
C13537 a_n232_53604# a_n232_53252# 0.0109f
C13538 AVDD a_14888_52548# 0.00166f
C13539 XA8.XA1.XA1.MN0.D a_19928_40228# 0.00155f
C13540 a_21080_40932# a_21080_40580# 0.0109f
C13541 a_9848_46564# a_9848_46212# 0.0109f
C13542 a_22448_46564# a_23600_46564# 0.00133f
C13543 XA8.XA3.MN0.G a_21080_46212# 0.155f
C13544 XA8.XA4.MN0.G a_21080_44804# 5.54e-19
C13545 XA1.XA4.MN0.G a_3440_44452# 0.00907f
C13546 XA7.XA1.XA5.MN2.G a_14888_41636# 0.128f
C13547 XA0.XA11.MN1.G a_11000_1742# 0.155f
C13548 XA3.XA4.MN0.D XA3.XA1.XA5.MN0.D 9.89e-19
C13549 VREF XA4.XA1.XA5.MP0.D 0.00202f
C13550 XA0.XA6.MP0.G a_920_42692# 5.5e-19
C13551 XA20.XA3a.MN0.D a_21080_45156# 3.15e-19
C13552 XA5.XA9.MN1.G XA6.XA9.MN1.G 0.0531f
C13553 XA1.XA10.MP0.G a_3440_51844# 5.59e-19
C13554 CK_SAMPLE a_n232_50436# 0.161f
C13555 AVDD XA4.XA6.MP0.G 5.98f
C13556 XB2.M1.G a_12368_686# 0.161f
C13557 XB1.M1.G CK_SAMPLE_BSSW 0.00269f
C13558 a_14960_1742# XB2.XA3.MN1.D 0.00685f
C13559 a_11000_1742# a_11000_1390# 0.0109f
C13560 XB1.XA0.MP0.D a_8408_1038# 0.081f
C13561 XB2.XA0.MP0.D a_14960_1390# 0.0749f
C13562 SARN XDAC2.X16ab.XRES16.B 55.3f
C13563 XA1.XA4.MN0.D XA1.XA1.XA1.MN0.D 0.00262f
C13564 XA20.XA3a.MN0.D XA1.XA1.XA4.MN0.D 1.1e-19
C13565 XA20.XA2a.MN0.D XA6.XA1.XA2.MP0.D 0.223f
C13566 a_16040_44804# a_17408_44804# 8.89e-19
C13567 a_3440_44804# a_3440_44452# 0.0109f
C13568 XA4.XA4.MN0.G a_11000_42340# 1.28e-19
C13569 D<8> a_n232_43044# 0.00321f
C13570 XA5.XA1.XA5.MN2.D a_13520_44100# 0.0893f
C13571 a_19928_45508# EN 3.34e-19
C13572 XA3.XA9.MN1.G a_7328_50084# 0.00281f
C13573 XA8.XA9.MN1.G XA8.XA6.MP0.D 0.0618f
C13574 AVDD a_16040_47268# 0.356f
C13575 XA0.XA10.MP0.G VREF 0.0134f
C13576 XA4.XA1.XA5.MN2.G XA3.XA6.MP2.D 0.00313f
C13577 XDAC1.X16ab.XRES2.B XDAC1.XC128b<2>.XRES2.B 1.67e-19
C13578 li_9184_23076# li_9184_22656# 0.00411f
C13579 XB1.XA4.MP0.D m3_n2104_3300# 0.0273f
C13580 a_19928_43748# a_19928_43396# 0.0109f
C13581 XA2.XA1.XA5.MN0.D a_5960_43396# 2.16e-19
C13582 XA2.XA1.XA5.MP0.D a_4808_43396# 2.16e-19
C13583 XA6.XA1.XA5.MN0.D XA6.XA1.XA5.MP0.D 0.00918f
C13584 XA20.XA2a.MN0.D XA4.XA1.XA1.MN0.D 0.0221f
C13585 EN XA5.XA1.XA4.MN1.D 3.17e-19
C13586 AVDD XA1.XA1.XA5.MN1.D 0.00889f
C13587 a_12368_50436# VREF 0.0035f
C13588 XA2.XA6.MP0.G a_5960_49732# 0.101f
C13589 XA2.XA6.MN0.D a_4808_49732# 0.00176f
C13590 XDAC1.XC1.XRES1B.B XDAC1.XC1.XRES1A.B 0.00438f
C13591 XDAC1.XC1.XRES4.B XDAC1.XC1.XRES16.B 0.0483f
C13592 XDAC1.XC1.XRES8.B XDAC1.XC1.XRES2.B 0.44f
C13593 XDAC2.XC1.XRES8.B li_14804_7512# 9.91e-20
C13594 XA3.XA3.MN0.G XDAC2.X16ab.XRES2.B 0.00405f
C13595 a_12368_43044# XA5.XA1.XA1.MN0.S 4.06e-20
C13596 XA2.XA1.XA2.MP0.D a_5960_40932# 4.25e-20
C13597 XA0.XA1.XA4.MP0.D a_920_41988# 0.00176f
C13598 XA5.XA1.XA4.MN0.D a_13520_42340# 0.0474f
C13599 a_920_42340# a_2288_42340# 8.89e-19
C13600 EN a_12368_40228# 0.0658f
C13601 D<0> a_19928_45860# 0.0675f
C13602 XA0.XA6.MP2.G XA0.XA1.XA5.MN2.D 0.0284f
C13603 a_7328_48676# a_7328_48324# 0.0109f
C13604 D<4> a_9848_45508# 0.0031f
C13605 XA7.XA1.XA5.MN2.G a_17408_45156# 7.1e-20
C13606 XA8.XA1.XA5.MN2.G a_16040_45156# 7.1e-20
C13607 XA20.XA9.MP0.D a_23600_43396# 0.00334f
C13608 AVDD a_16040_41636# 0.404f
C13609 XA7.XA6.MP0.G XA2.XA3.MN0.G 0.0653f
C13610 VREF a_13520_47620# 7.12e-19
C13611 AVDD a_920_53252# 0.364f
C13612 CK_SAMPLE XA20.XA10.MN0.D 0.00225f
C13613 a_22448_53956# a_23600_53956# 0.00133f
C13614 a_9848_53956# XA4.XA12.MP0.G 0.0704f
C13615 a_11000_53956# XA5.XA11.MN1.G 0.0442f
C13616 XA0.XA1.XA1.MN0.D a_920_40932# 8.29e-20
C13617 SARP XDAC1.XC32a<0>.XRES16.B 55.3f
C13618 XA7.XA6.MP0.G a_17408_43748# 5.5e-19
C13619 D<5> XA3.XA1.XA4.MP1.D 7.43e-19
C13620 VREF a_2288_44100# 0.0251f
C13621 XA1.XA4.MN0.G a_3440_45508# 0.0104f
C13622 XA8.XA4.MN0.G a_19928_45860# 0.0146f
C13623 AVDD a_9560_686# 0.00165f
C13624 XA8.XA7.MP0.G a_22448_42692# 0.00119f
C13625 a_19928_47268# XA8.XA3.MN0.G 2.69e-19
C13626 a_3440_46916# XA1.XA3.MN0.G 0.0666f
C13627 XA3.XA1.XA5.MN2.G XA2.XA1.XA4.MN0.D 7.2e-19
C13628 D<1> a_17408_43044# 7.77e-20
C13629 XA20.XA10.MN1.D a_23600_39876# 7.39e-19
C13630 XA2.XA1.XA5.MN2.G XA2.XA1.XA4.MP0.D 6.33e-19
C13631 XA0.XA10.MP0.G a_920_52548# 0.07f
C13632 XA5.XA10.MP0.G XA6.XA10.MP0.G 0.00217f
C13633 AVDD XA2.XA6.MP2.D 0.172f
C13634 CK_SAMPLE XA6.XA1.XA5.MN2.G 0.0595f
C13635 a_9560_3502# XB1.M1.G 5.7e-19
C13636 a_8408_3502# XB1.XA4.MP0.D 0.00426f
C13637 a_12368_2798# a_13808_2798# 8e-19
C13638 a_9560_2798# XB1.XA1.MP0.D 0.0153f
C13639 a_8408_2798# XB1.XA1.MN0.D 0.0674f
C13640 a_14960_3502# XB2.XA1.MP0.D 1.47e-19
C13641 XA2.XA1.XA5.MN2.D a_5960_45156# 0.155f
C13642 XA6.XA4.MN0.G a_16040_43044# 0.0222f
C13643 XA8.XA1.XA5.MN2.G a_19928_39876# 0.00169f
C13644 XA5.XA6.MP0.G a_12368_41284# 4.24e-19
C13645 XA20.XA3a.MN0.D a_12368_43396# 0.00213f
C13646 a_16040_51844# XA7.XA1.XA5.MN2.G 8.87e-19
C13647 XA6.XA7.MP0.D a_16040_51140# 0.00224f
C13648 CK_SAMPLE a_n232_48676# 4.46e-19
C13649 AVDD a_14888_48324# 0.00131f
C13650 a_5960_51492# a_7328_51492# 8.89e-19
C13651 XA6.XA8.MP0.D a_16040_51492# 0.00224f
C13652 a_11000_53604# VREF 0.00351f
C13653 XA20.XA3a.MN0.D a_11000_40932# 0.0658f
C13654 XA4.XA1.XA5.MN2.D a_11000_42692# 7.44e-20
C13655 XA20.XA2a.MN0.D a_18560_41988# 0.0861f
C13656 XA6.XA1.XA5.MP1.D a_16040_43748# 0.049f
C13657 XA2.XA3.MN0.G XA1.XA1.XA1.MN0.S 0.00103f
C13658 EN XA2.XA1.XA5.MN0.D 0.0063f
C13659 XA1.XA1.XA5.MN1.D XA1.XA1.XA2.MP0.D 0.0102f
C13660 XA1.XA1.XA5.MP1.D XA1.XA1.XA5.MP0.D 0.0488f
C13661 a_18560_50436# a_19928_50436# 8.89e-19
C13662 a_4808_50436# XA2.XA6.MN0.D 0.00176f
C13663 a_5960_50436# XA2.XA6.MP0.G 0.0662f
C13664 a_16040_50788# XA6.XA6.MP0.G 1.34e-19
C13665 AVDD a_18560_45156# 0.00125f
C13666 a_7328_51140# VREF 0.00383f
C13667 XA7.XA1.XA4.MP1.D a_17408_42692# 0.049f
C13668 XA7.XA1.XA2.MP0.D a_18560_41988# 0.0568f
C13669 XA3.XA1.XA2.MP0.D a_8480_41636# 0.00316f
C13670 XA2.XA1.XA4.MN1.D XA2.XA1.XA4.MN0.D 0.0488f
C13671 EN a_21080_41284# 0.00558f
C13672 AVDD XA0.XA1.XA4.MP0.D 0.152f
C13673 XA3.XA4.MN0.D a_8480_48676# 0.158f
C13674 VREF a_12368_48676# 0.0191f
C13675 D<2> XA1.XA3.MN0.G 0.0258f
C13676 a_n232_49028# a_920_49028# 0.00133f
C13677 D<6> a_4808_46564# 0.0551f
C13678 AVDD CK_SAMPLE 5.8f
C13679 a_16040_41636# a_16040_41284# 0.0109f
C13680 XA8.XA4.MN0.G a_18560_46916# 2.84e-19
C13681 XA7.XA4.MN0.G a_19928_46916# 2.84e-19
C13682 XA2.XA4.MN0.G XA1.XA3.MN0.G 0.00444f
C13683 XA1.XA4.MN0.G XA2.XA3.MN0.G 0.00499f
C13684 a_19928_47620# a_21080_47620# 0.00133f
C13685 XA5.XA1.XA5.MN2.G a_11000_43396# 0.00442f
C13686 VREF XA2.XA1.XA5.MN2.D 0.341f
C13687 XA1.XA4.MN0.D XA1.XA1.XA5.MN2.D 0.0264f
C13688 AVDD a_22448_39876# 0.438f
C13689 D<2> a_16040_43748# 7.76e-20
C13690 XA6.XA11.MP0.D a_16040_52900# 0.00176f
C13691 a_5960_53252# a_5960_52900# 0.0109f
C13692 XA8.XA11.MN1.G a_18560_52548# 9.76e-19
C13693 AVDD a_17408_51844# 0.387f
C13694 XA0.XA11.MN1.G XA0.XA10.MP0.G 7.66e-19
C13695 XA2.XA12.MP0.G XA2.XA9.MN1.G 4.5e-19
C13696 a_14888_40228# a_14888_39876# 0.0109f
C13697 XA0.XA4.MN0.D a_n232_42692# 9.25e-20
C13698 XA20.XA2a.MN0.D XA6.XA1.XA5.MN2.D 8.92e-20
C13699 a_14888_45860# a_16040_45860# 0.00133f
C13700 XA5.XA4.MN0.G a_12368_43748# 6.3e-19
C13701 XA20.XA3a.MN0.D XA2.XA1.XA5.MN1.D 2.15e-19
C13702 XA1.XA3.MN0.G a_4808_44804# 4.4e-20
C13703 XA2.XA3.MN0.G a_3440_44804# 2.51e-19
C13704 XA5.XA1.XA5.MN2.G a_9848_40932# 6.44e-19
C13705 XA4.XA1.XA5.MN2.G a_11000_40932# 1.69e-19
C13706 D<4> a_11000_41284# 7.76e-20
C13707 AVDD a_920_49380# 0.356f
C13708 DONE VREF 0.108f
C13709 XA4.XA9.MN1.G a_9848_51492# 0.0118f
C13710 XA20.XA2.MN1.D a_22448_43748# 0.00253f
C13711 XA20.XA2a.MN0.D a_3440_42692# 0.00563f
C13712 XA0.XA1.XA5.MN2.D a_n232_43396# 1.28e-19
C13713 XA0.XA6.MP2.G XDAC1.XC64b<1>.XRES4.B 4.06e-21
C13714 SARN li_14804_13860# 0.00103f
C13715 a_8480_44100# a_9848_44100# 8.89e-19
C13716 a_18560_44452# EN 0.00154f
C13717 AVDD a_16040_46212# 0.356f
C13718 XA5.XA1.XA5.MN2.G XA4.XA6.MP0.G 0.0959f
C13719 XA1.XA7.MP0.D VREF 0.0234f
C13720 XDAC2.XC128a<1>.XRES8.B XDAC2.XC128a<1>.XRES2.B 0.44f
C13721 XDAC2.XC128a<1>.XRES4.B XDAC2.XC128a<1>.XRES16.B 0.0483f
C13722 XDAC2.XC128a<1>.XRES1B.B XDAC2.XC128a<1>.XRES1A.B 0.00438f
C13723 XA20.XA2a.MN0.D a_n232_39876# 1.09e-19
C13724 a_8480_43044# a_9848_43044# 8.89e-19
C13725 XA0.XA6.MP0.G XDAC2.XC1.XRES4.B 0.00405f
C13726 EN a_4808_41988# 1.25e-19
C13727 XA6.XA6.MP0.G a_16040_49028# 0.0307f
C13728 D<5> XA20.XA3a.MN0.D 0.0703f
C13729 AVDD a_9848_43396# 0.00125f
C13730 XA2.XA6.MP0.G a_5960_48676# 0.0881f
C13731 a_n232_49732# a_n232_49380# 0.0109f
C13732 a_7328_49732# XA3.XA4.MN0.D 0.0674f
C13733 a_11000_49732# VREF 0.029f
C13734 a_19928_41988# a_21080_41988# 0.00133f
C13735 AVDD a_8480_40932# 0.00125f
C13736 XA3.XA1.XA5.MN2.G XA2.XA1.XA5.MP1.D 0.00329f
C13737 XA8.XA7.MP0.G EN 0.793f
C13738 XA4.XA4.MN0.G a_11000_47972# 0.155f
C13739 XA4.XA4.MN0.D a_9848_46564# 4.06e-19
C13740 VREF a_14888_46564# 7.39e-19
C13741 XA4.XA12.MP0.G a_11000_53252# 0.00276f
C13742 XA5.XA11.MN1.G a_12368_53252# 0.0762f
C13743 a_17408_53604# a_18560_53604# 0.00133f
C13744 AVDD a_13520_52548# 0.00166f
C13745 a_7328_40580# a_8480_40580# 0.00133f
C13746 XA8.XA3.MN0.G a_19928_46212# 0.157f
C13747 XA1.XA3.MN0.G a_3440_45860# 0.162f
C13748 XA1.XA4.MN0.G a_2288_44452# 5.54e-19
C13749 XA8.XA4.MN0.G a_19928_44804# 0.00858f
C13750 XA6.XA1.XA5.MN2.G a_14888_41636# 0.00417f
C13751 XA0.XA11.MN1.G a_9560_1742# 0.00212f
C13752 XA3.XA4.MN0.D XA3.XA1.XA5.MP0.D 9.71e-19
C13753 XA0.XA6.MP0.G a_n232_42692# 7.76e-20
C13754 SARN a_23600_40932# 5.16e-19
C13755 XA1.XA10.MP0.G a_2288_51844# 0.00224f
C13756 XA6.XA10.MP0.G XA6.XA7.MP0.D 0.0601f
C13757 AVDD XA3.XA6.MN0.D 3.13e-19
C13758 XA5.XA9.MN1.G XA5.XA9.MN0.D 0.034f
C13759 a_13520_52548# a_13520_52196# 0.0109f
C13760 SAR_IP a_11000_n18# 0.0347f
C13761 XB1.XA3.MN0.S XB1.XA3.MN1.D 0.0944f
C13762 a_13808_1742# XB2.XA3.MN1.D 0.00176f
C13763 XB2.XA0.MP0.D a_13808_1390# 0.0735f
C13764 XA20.XA3a.MN0.D XA1.XA1.XA4.MP0.D 1.1e-19
C13765 XA4.XA4.MN0.G a_9848_42340# 7.97e-19
C13766 XA5.XA1.XA5.MN2.D a_12368_44100# 0.124f
C13767 a_18560_45508# EN 3.34e-19
C13768 XA7.XA7.MP0.D a_18560_50436# 1.37e-19
C13769 XA8.XA9.MN1.G XA8.XA6.MN0.D 0.0615f
C13770 a_920_51140# XA0.XA6.MP2.D 0.00176f
C13771 a_13520_51140# a_14888_51140# 8.89e-19
C13772 AVDD a_14888_47268# 0.00125f
C13773 XA4.XA1.XA5.MN2.G D<5> 0.691f
C13774 XB1.XA4.MP0.D m3_7544_3476# 0.106f
C13775 XA2.XA1.XA5.MN0.D a_4808_43396# 0.0474f
C13776 XA6.XA1.XA2.MP0.D XA6.XA1.XA5.MP0.D 4.34e-19
C13777 XA20.XA2a.MN0.D XA3.XA1.XA1.MN0.D 0.022f
C13778 EN XA5.XA1.XA4.MP1.D 0.0386f
C13779 XA6.XA6.MN0.D a_14888_50084# 0.0488f
C13780 XA6.XA6.MP0.G a_16040_50084# 0.159f
C13781 AVDD XA1.XA1.XA5.MP1.D 0.0889f
C13782 a_n232_50084# a_920_50084# 0.00133f
C13783 a_11000_50436# VREF 0.0035f
C13784 XA2.XA6.MP0.G a_4808_49732# 0.00239f
C13785 D<8> li_14804_24300# 3.5e-20
C13786 XA5.XA1.XA4.MN0.D a_12368_42340# 2.16e-19
C13787 XA5.XA1.XA4.MP0.D a_13520_42340# 2.16e-19
C13788 EN a_11000_40228# 0.0674f
C13789 D<0> a_18560_45860# 1.06e-19
C13790 XA7.XA1.XA5.MN2.G a_16040_45156# 0.00486f
C13791 a_18560_48676# a_19928_48676# 8.89e-19
C13792 XA20.XA9.MP0.D a_22448_43396# 0.0736f
C13793 AVDD a_14888_41636# 0.00125f
C13794 XA7.XA6.MP0.G XA1.XA3.MN0.G 0.0302f
C13795 VREF a_12368_47620# 0.0671f
C13796 XA3.XA4.MN0.D a_8480_47620# 0.0396f
C13797 AVDD a_n232_53252# 0.00154f
C13798 CK_SAMPLE XA20.XA10.MN1.D 0.0445f
C13799 a_9848_53956# XA5.XA11.MN1.G 0.0224f
C13800 a_12368_41284# a_12368_40932# 0.0109f
C13801 XA0.XA1.XA1.MN0.D a_n232_40932# 0.0535f
C13802 VREF a_920_44100# 0.0251f
C13803 XA2.XA6.MP0.G XA2.XA1.XA5.MP0.D 0.00121f
C13804 XA1.XA4.MN0.G a_2288_45508# 6.57e-19
C13805 XA7.XA4.MN0.G a_19928_45860# 2.2e-19
C13806 XA8.XA4.MN0.G a_18560_45860# 2.2e-19
C13807 AVDD a_8408_686# 0.37f
C13808 XA8.XA7.MP0.G a_21080_42692# 0.00442f
C13809 a_13520_46916# a_14888_46916# 8.89e-19
C13810 a_2288_46916# XA1.XA3.MN0.G 0.0674f
C13811 XA2.XA1.XA5.MN2.G XA2.XA1.XA4.MN0.D 0.00313f
C13812 DONE a_21080_51140# 9.73e-19
C13813 a_12368_52900# a_12368_52548# 0.0109f
C13814 XA0.XA10.MP0.G a_n232_52548# 0.128f
C13815 a_n232_52900# XA0.XA9.MN1.G 0.00113f
C13816 AVDD XA2.XA6.MN2.D 3.77e-19
C13817 CK_SAMPLE XA5.XA1.XA5.MN2.G 0.0595f
C13818 a_8408_2798# XB1.XA1.MP0.D 0.0317f
C13819 XB2.XA2.MN0.G XB2.XA1.MN0.D 0.0103f
C13820 a_13808_3502# XB2.XA1.MP0.D 2.12e-19
C13821 a_16040_45508# a_16040_45156# 0.0109f
C13822 XA2.XA1.XA5.MN2.D a_4808_45156# 0.153f
C13823 XA7.XA1.XA5.MN2.D XA8.XA1.XA5.MN2.D 0.00869f
C13824 XA6.XA4.MN0.G a_14888_43044# 0.0409f
C13825 XA8.XA1.XA5.MN2.G a_18560_39876# 2.97e-20
C13826 XA3.XA4.MN0.D a_8480_41988# 9.24e-20
C13827 XA20.XA3a.MN0.D a_11000_43396# 0.00213f
C13828 XA7.XA9.MN1.G XA7.XA6.MN2.D 0.126f
C13829 XA6.XA7.MP0.D a_14888_51140# 0.00388f
C13830 AVDD a_13520_48324# 0.00131f
C13831 a_23600_51844# a_23600_51492# 0.0109f
C13832 XA6.XA8.MP0.D a_14888_51492# 0.00224f
C13833 XDAC1.XC64b<1>.XRES1B.B XDAC1.X16ab.XRES1B.B 0.00444f
C13834 XDAC1.XC64b<1>.XRES4.B XDAC1.XC64b<1>.XRES1A.B 0.0197f
C13835 li_9184_28392# li_9184_27780# 0.00271f
C13836 XDAC1.XC64b<1>.XRES8.B XDAC1.XC64b<1>.XRES16.B 0.0904f
C13837 XA20.XA3a.MN0.D a_9848_40932# 0.0739f
C13838 XA20.XA2a.MN0.D a_17408_41988# 0.00302f
C13839 XA6.XA1.XA5.MP1.D a_14888_43748# 2.16e-19
C13840 XA6.XA1.XA5.MN1.D a_16040_43748# 2.16e-19
C13841 a_3440_43748# a_4808_43748# 8.89e-19
C13842 XA0.XA6.MP2.G li_9184_19176# 0.00508f
C13843 XA1.XA3.MN0.G XA1.XA1.XA1.MN0.S 0.00995f
C13844 a_13520_44100# XA5.XA1.XA2.MP0.D 2.92e-19
C13845 XA1.XA1.XA5.MP1.D XA1.XA1.XA2.MP0.D 6.52e-20
C13846 EN XA2.XA1.XA2.MP0.D 0.03f
C13847 a_4808_50436# XA2.XA6.MP0.G 3.02e-20
C13848 a_14888_50788# XA6.XA6.MP0.G 1.75e-20
C13849 AVDD a_17408_45156# 0.356f
C13850 a_5960_51140# VREF 0.00383f
C13851 D<7> a_3440_49732# 7.01e-19
C13852 XA8.XA1.XA5.MN2.G XA7.XA4.MN0.D 0.0939f
C13853 a_4808_42692# a_5960_42692# 0.00133f
C13854 XA7.XA1.XA2.MP0.D a_17408_41988# 0.0219f
C13855 XA3.XA1.XA2.MP0.D a_7328_41636# 0.00224f
C13856 SARP a_23600_40932# 0.159f
C13857 XA0.XA4.MN0.D XDAC1.XC1.XRES4.B 0.00405f
C13858 XA3.XA4.MN0.D a_7328_48676# 0.154f
C13859 VREF a_11000_48676# 0.0191f
C13860 AVDD XA0.XA1.XA4.MN0.D 0.00889f
C13861 D<2> D<8> 0.0322f
C13862 XA2.XA6.MP0.G a_5960_47620# 6.35e-19
C13863 D<3> XA3.XA3.MN0.G 0.12f
C13864 XA4.XA6.MP0.G XA20.XA3a.MN0.D 0.0771f
C13865 a_12368_49380# a_12368_49028# 0.0109f
C13866 AVDD a_23600_54308# 0.00154f
C13867 a_3440_54308# a_4808_54308# 8.89e-19
C13868 SARP XDAC1.X16ab.XRES16.B 55.3f
C13869 XA1.XA1.XA1.MP2.D a_2288_41284# 0.0465f
C13870 XA1.XA1.XA1.MN0.S a_3440_41284# 0.0674f
C13871 XA5.XA1.XA5.MN2.G a_9848_43396# 1.95e-19
C13872 a_7328_47620# a_7328_47268# 0.0109f
C13873 XA1.XA4.MN0.G XA1.XA3.MN0.G 0.639f
C13874 XA7.XA4.MN0.G a_18560_46916# 0.0885f
C13875 VREF XA1.XA1.XA5.MN2.D 0.341f
C13876 AVDD a_21080_39876# 0.44f
C13877 D<2> a_14888_43748# 6.49e-19
C13878 a_16040_53252# XA6.XA10.MP0.D 0.0661f
C13879 XA8.XA11.MN1.G a_17408_52548# 7.25e-20
C13880 AVDD a_16040_51844# 0.387f
C13881 XA3.XA11.MN1.G XA2.XA9.MN1.G 0.00116f
C13882 a_920_39876# a_2288_39876# 8.89e-19
C13883 XA2.XA6.MP0.G a_5960_41988# 5.5e-19
C13884 SARN a_13808_3502# 0.00116f
C13885 XA20.XA2a.MN0.D XA5.XA1.XA5.MN2.D 8.92e-20
C13886 a_2288_45860# a_2288_45508# 0.0109f
C13887 XA6.XA6.MP0.G a_16040_42340# 5.5e-19
C13888 XA1.XA3.MN0.G a_3440_44804# 0.0433f
C13889 XA8.XA3.MN0.G a_21080_45156# 0.0546f
C13890 XA20.XA3a.MN0.D XA1.XA1.XA5.MN1.D 2.15e-19
C13891 XA0.XA6.MP2.G XA0.XA1.XA1.MN0.D 0.0192f
C13892 XA4.XA1.XA5.MN2.G a_9848_40932# 0.00729f
C13893 D<4> a_9848_41284# 6.49e-19
C13894 AVDD a_n232_49380# 0.00159f
C13895 XA20.XA11.MN0.D VREF 0.00269f
C13896 a_14888_52196# a_14888_51844# 0.0109f
C13897 a_3440_52196# XA1.XA8.MP0.D 2.11e-19
C13898 XA4.XA9.MN1.G a_8480_51492# 2.84e-19
C13899 a_12368_52548# XA6.XA1.XA5.MN2.G 1.75e-19
C13900 XA1.XA7.MP0.D a_3440_51844# 0.159f
C13901 XA6.XA7.MP0.D XA7.XA7.MP0.D 0.00435f
C13902 XA20.XA2a.MN0.D a_2288_42692# 0.00457f
C13903 D<7> XDAC1.XC64b<1>.XRES1B.B 0.00405f
C13904 a_21080_44452# a_21080_44100# 0.0109f
C13905 a_17408_44452# EN 0.00173f
C13906 AVDD a_14888_46212# 0.00125f
C13907 XA4.XA1.XA5.MN2.G XA4.XA6.MP0.G 0.00254f
C13908 a_17408_51492# XA7.XA6.MP0.G 4.06e-20
C13909 XA0.XA7.MP0.D VREF 0.0234f
C13910 XA1.XA6.MP2.D a_2288_50436# 0.00176f
C13911 D<7> a_3440_50436# 5.7e-19
C13912 XA5.XA6.MP2.D a_12368_50788# 0.049f
C13913 XA8.XA1.XA2.MP0.D XA8.XA1.XA4.MP1.D 4.34e-19
C13914 a_21080_43396# a_21080_43044# 0.0109f
C13915 EN a_3440_41988# 1.25e-19
C13916 XA6.XA6.MP0.G a_14888_49028# 0.0137f
C13917 AVDD a_8480_43396# 0.00125f
C13918 XA2.XA6.MP0.G a_4808_48676# 0.0651f
C13919 a_17408_49732# a_18560_49732# 0.00133f
C13920 a_7328_41988# a_7328_41636# 0.0109f
C13921 a_7328_42340# XA3.XA1.XA1.MN0.S 1.34e-19
C13922 AVDD a_7328_40932# 0.358f
C13923 XA2.XA1.XA5.MN2.G XA2.XA1.XA5.MP1.D 5.21e-20
C13924 SARN a_23600_43396# 0.0017f
C13925 XA3.XA1.XA5.MN2.G XA2.XA1.XA5.MN1.D 6.68e-19
C13926 XA8.XA1.XA5.MN2.G EN 0.898f
C13927 a_920_47972# a_2288_47972# 8.89e-19
C13928 XA4.XA4.MN0.G a_9848_47972# 0.153f
C13929 a_19928_48324# a_19928_47972# 0.0109f
C13930 VREF a_13520_46564# 7.39e-19
C13931 a_5960_53604# XA2.XA11.MP0.D 0.00176f
C13932 XA5.XA11.MN1.G a_11000_53252# 0.00648f
C13933 XA4.XA12.MP0.G a_9848_53252# 0.0661f
C13934 AVDD a_12368_52548# 0.405f
C13935 XA7.XA1.XA1.MN0.D a_18560_40228# 0.00155f
C13936 a_19928_40932# a_19928_40580# 0.0109f
C13937 XA6.XA1.XA5.MN2.G a_13520_41636# 0.131f
C13938 XA1.XA3.MN0.G a_2288_45860# 0.155f
C13939 XA8.XA4.MN0.G a_18560_44804# 2.2e-19
C13940 XA7.XA4.MN0.G a_19928_44804# 2.2e-19
C13941 XA3.XA4.MN0.D XA3.XA1.XA2.MP0.D 0.0111f
C13942 a_21080_46564# a_22448_46564# 8.89e-19
C13943 a_8480_46564# a_8480_46212# 0.0109f
C13944 AVDD XA3.XA6.MP0.D 0.144f
C13945 CK_SAMPLE a_22448_50788# 0.00273f
C13946 XA0.XA9.MN1.G a_920_52196# 0.0681f
C13947 XA0.XA9.MN0.D a_n232_52196# 0.0492f
C13948 XB2.XA4.MP0.D a_14960_1038# 0.00161f
C13949 a_13808_1742# XB2.XA3.MN0.S 0.0703f
C13950 a_9560_1742# a_9560_1390# 0.0109f
C13951 XA20.XA3a.MN0.D XA0.XA1.XA4.MP0.D 1.1e-19
C13952 a_14888_44804# a_16040_44804# 0.00133f
C13953 a_2288_44804# a_2288_44452# 0.0109f
C13954 XA3.XA6.MP0.G a_8480_40228# 3.45e-20
C13955 XA6.XA3.MN0.G a_14888_43396# 6.8e-20
C13956 a_17408_45508# EN 1.42e-19
C13957 XA7.XA6.MP0.G a_18560_40580# 7.76e-20
C13958 SARN li_14804_24300# 0.00103f
C13959 a_16040_51492# D<2> 2.41e-19
C13960 XA8.XA9.MN1.G XA8.XA6.MP0.G 0.0725f
C13961 AVDD a_13520_47268# 0.00125f
C13962 a_22448_52900# VREF 0.00125f
C13963 XA3.XA1.XA5.MN2.G D<5> 0.0713f
C13964 XB1.XA4.MP0.D m3_7472_3476# 0.0634f
C13965 XDAC2.X16ab.XRES1A.B XDAC2.XC128b<2>.XRES1B.B 0.617f
C13966 a_18560_43748# a_18560_43396# 0.0109f
C13967 XA2.XA1.XA2.MP0.D a_4808_43396# 0.0945f
C13968 XA6.XA1.XA2.MP0.D XA6.XA1.XA5.MN0.D 0.056f
C13969 XA20.XA2a.MN0.D XA3.XA1.XA1.MP1.D 0.00946f
C13970 EN XA4.XA1.XA4.MP1.D 0.0386f
C13971 XA6.XA6.MP0.G a_14888_50084# 6.4e-20
C13972 AVDD XA0.XA1.XA5.MP1.D 0.0889f
C13973 D<3> a_13520_49028# 5.7e-19
C13974 D<7> a_3440_48676# 3.48e-19
C13975 XA6.XA1.XA5.MN2.G a_12368_48324# 0.00455f
C13976 XDAC2.XC1.XRES4.B XDAC2.XC1.XRES2.B 0.0307f
C13977 li_14804_8124# li_14804_7512# 0.00271f
C13978 XDAC2.XC64a<0>.XRES1A.B XDAC2.XC1.XRES1A.B 0.00444f
C13979 XDAC2.XC1.XRES1B.B XDAC2.XC1.XRES16.B 0.0381f
C13980 XDAC1.XC1.XRES8.B li_9184_7512# 9.91e-20
C13981 XA0.XA1.XA4.MN0.D a_n232_41988# 0.00176f
C13982 XA5.XA1.XA4.MP0.D a_12368_42340# 0.049f
C13983 a_n232_42340# a_920_42340# 0.00133f
C13984 XA7.XA1.XA5.MN2.G a_14888_45156# 1.95e-19
C13985 a_5960_48676# a_5960_48324# 0.0109f
C13986 XA6.XA6.MP0.G XA3.XA3.MN0.G 0.0337f
C13987 XA20.XA9.MP0.D a_21080_43396# 5.7e-20
C13988 AVDD a_13520_41636# 0.00125f
C13989 XA7.XA6.MP0.G D<8> 0.132f
C13990 VREF a_11000_47620# 0.0671f
C13991 XA3.XA4.MN0.D a_7328_47620# 0.00498f
C13992 DONE a_23600_53604# 1.69e-19
C13993 AVDD XA8.XA11.MP0.D 0.19f
C13994 a_23600_54308# XA20.XA10.MN1.D 7.49e-19
C13995 CK_SAMPLE XA8.XA12.MP0.G 0.00163f
C13996 a_21080_53956# a_22448_53956# 8.89e-19
C13997 XA4.XA1.XA1.MN0.S a_11000_40580# 0.0318f
C13998 SARP li_9184_13860# 0.00103f
C13999 XA0.XA4.MN0.D a_920_44100# 9.14e-20
C14000 XA2.XA6.MP0.G XA2.XA1.XA5.MN0.D 7.41e-19
C14001 XA7.XA4.MN0.G a_18560_45860# 0.0146f
C14002 AVDD a_14960_1038# 0.489f
C14003 XA8.XA7.MP0.G a_19928_42692# 1.95e-19
C14004 a_18560_47268# XA7.XA3.MN0.G 2.69e-19
C14005 XA8.XA1.XA5.MN2.G a_21080_42692# 1.97e-19
C14006 XA2.XA1.XA5.MN2.G XA1.XA1.XA4.MN0.D 7.72e-19
C14007 XA3.XA10.MP0.D XA3.XA9.MN1.G 0.00406f
C14008 DONE a_19928_51140# 3.16e-19
C14009 XA4.XA10.MP0.G XA5.XA10.MP0.G 0.00217f
C14010 a_18560_53252# XA7.XA9.MN1.G 5.25e-19
C14011 AVDD D<6> 2.23f
C14012 CK_SAMPLE XA4.XA1.XA5.MN2.G 0.0595f
C14013 a_9560_3854# XB1.M1.G 3.5e-19
C14014 a_8408_3854# XB1.XA4.MP0.D 0.0036f
C14015 a_11000_2798# a_12368_2798# 8.89e-19
C14016 a_14960_3854# XB2.XA1.MP0.D 7.02e-20
C14017 XA7.XA1.XA5.MN2.G a_18560_39876# 0.00325f
C14018 XA8.XA1.XA5.MN2.G a_17408_39876# 8.8e-19
C14019 XA3.XA4.MN0.D a_7328_41988# 9.15e-20
C14020 SARN a_13808_334# 2.97e-20
C14021 XA20.XA3a.MN0.D a_9848_43396# 0.0736f
C14022 a_4808_51492# a_5960_51492# 0.00133f
C14023 XA7.XA9.MN1.G XA7.XA6.MP2.D 0.0618f
C14024 AVDD a_12368_48324# 0.359f
C14025 XA2.XA9.MN1.G a_5960_50788# 0.00281f
C14026 SARN D<2> 0.027f
C14027 XA20.XA3a.MN0.D a_8480_40932# 0.0723f
C14028 XA20.XA2a.MN0.D a_16040_41988# 0.00302f
C14029 SARP a_23600_43396# 0.158f
C14030 XA6.XA1.XA5.MN1.D a_14888_43748# 0.0494f
C14031 EN XA1.XA1.XA5.MN0.D 0.0063f
C14032 m3_26048_132# AVSS 0.00417f
C14033 m3_25976_132# AVSS 0.00167f $ **FLOATING
C14034 m3_16544_308# AVSS 0.00167f $ **FLOATING
C14035 m3_16472_308# AVSS 0.0025f
C14036 m3_26048_1188# AVSS 0.00417f
C14037 m3_25976_1188# AVSS 0.00167f $ **FLOATING
C14038 m3_16544_1364# AVSS 0.00167f $ **FLOATING
C14039 m3_16472_1364# AVSS 0.0025f
C14040 m3_26048_2244# AVSS 0.00417f
C14041 m3_25976_2244# AVSS 0.00167f $ **FLOATING
C14042 m3_16544_2420# AVSS 0.00167f $ **FLOATING
C14043 m3_16472_2420# AVSS 0.0025f
C14044 m3_26048_3300# AVSS 0.00417f
C14045 m3_25976_3300# AVSS 0.00167f $ **FLOATING
C14046 m3_16544_3476# AVSS 0.00167f $ **FLOATING
C14047 m3_16472_3476# AVSS 0.0025f
C14048 m3_26048_4356# AVSS 0.00417f
C14049 m3_25976_4356# AVSS 0.00167f $ **FLOATING
C14050 m3_16544_4532# AVSS 0.00187f $ **FLOATING
C14051 m3_16472_4532# AVSS 0.00271f
C14052 m3_n1960_132# AVSS 0.00167f $ **FLOATING
C14053 m3_n2104_132# AVSS 0.00417f
C14054 m3_7544_308# AVSS 0.0025f
C14055 m3_7472_308# AVSS 0.00167f $ **FLOATING
C14056 m3_n1960_1188# AVSS 0.00167f $ **FLOATING
C14057 m3_n2104_1188# AVSS 0.00417f
C14058 m3_7544_1364# AVSS 0.0025f
C14059 m3_7472_1364# AVSS 0.00167f $ **FLOATING
C14060 m3_n1960_2244# AVSS 0.00167f $ **FLOATING
C14061 m3_n2104_2244# AVSS 0.00417f
C14062 m3_7544_2420# AVSS 0.0025f
C14063 m3_7472_2420# AVSS 0.00167f $ **FLOATING
C14064 m3_n1960_3300# AVSS 0.00167f $ **FLOATING
C14065 m3_n2104_3300# AVSS 0.00417f
C14066 m3_7544_3476# AVSS 0.0025f
C14067 m3_7472_3476# AVSS 0.00167f $ **FLOATING
C14068 m3_n1960_4356# AVSS 0.00167f $ **FLOATING
C14069 m3_n2104_4356# AVSS 0.00417f
C14070 m3_7544_4532# AVSS 0.00271f
C14071 m3_7472_4532# AVSS 0.00187f $ **FLOATING
C14072 li_14804_5676# AVSS 0.0349f $ **FLOATING
C14073 li_9184_5676# AVSS 0.0349f $ **FLOATING
C14074 XDAC2.XC1.XRES1A.B AVSS 8.27f
C14075 XDAC1.XC1.XRES1A.B AVSS 8.27f
C14076 li_14804_6288# AVSS 0.0311f $ **FLOATING
C14077 li_9184_6288# AVSS 0.0311f $ **FLOATING
C14078 XDAC2.XC1.XRES16.B AVSS 22.8f
C14079 XDAC1.XC1.XRES16.B AVSS 22.8f
C14080 li_14804_6900# AVSS 0.031f $ **FLOATING
C14081 li_9184_6900# AVSS 0.031f $ **FLOATING
C14082 XDAC2.XC1.XRES2.B AVSS 9.09f
C14083 XDAC1.XC1.XRES2.B AVSS 9.09f
C14084 li_14804_7512# AVSS 0.031f $ **FLOATING
C14085 li_9184_7512# AVSS 0.031f $ **FLOATING
C14086 XDAC2.XC1.XRES8.B AVSS 15f
C14087 XDAC1.XC1.XRES8.B AVSS 15f
C14088 li_14804_8124# AVSS 0.0311f $ **FLOATING
C14089 li_9184_8124# AVSS 0.0311f $ **FLOATING
C14090 XDAC2.XC1.XRES4.B AVSS 11.1f
C14091 XDAC1.XC1.XRES4.B AVSS 11.1f
C14092 li_14804_8736# AVSS 0.0299f $ **FLOATING
C14093 li_9184_8736# AVSS 0.0299f $ **FLOATING
C14094 XDAC2.XC1.XRES1B.B AVSS 8.07f
C14095 XDAC1.XC1.XRES1B.B AVSS 8.07f
C14096 li_14804_9156# AVSS 0.0299f $ **FLOATING
C14097 li_9184_9156# AVSS 0.0299f $ **FLOATING
C14098 XDAC2.XC64a<0>.XRES1A.B AVSS 8.06f
C14099 XDAC1.XC64a<0>.XRES1A.B AVSS 8.06f
C14100 li_14804_9768# AVSS 0.0311f $ **FLOATING
C14101 li_9184_9768# AVSS 0.0311f $ **FLOATING
C14102 XDAC2.XC64a<0>.XRES16.B AVSS 22.8f
C14103 XDAC1.XC64a<0>.XRES16.B AVSS 22.8f
C14104 li_14804_10380# AVSS 0.031f $ **FLOATING
C14105 li_9184_10380# AVSS 0.031f $ **FLOATING
C14106 XDAC2.XC64a<0>.XRES2.B AVSS 9.09f
C14107 XDAC1.XC64a<0>.XRES2.B AVSS 9.09f
C14108 li_14804_10992# AVSS 0.031f $ **FLOATING
C14109 li_9184_10992# AVSS 0.031f $ **FLOATING
C14110 XDAC2.XC64a<0>.XRES8.B AVSS 15f
C14111 XDAC1.XC64a<0>.XRES8.B AVSS 15f
C14112 li_14804_11604# AVSS 0.0311f $ **FLOATING
C14113 li_9184_11604# AVSS 0.0311f $ **FLOATING
C14114 XDAC2.XC64a<0>.XRES4.B AVSS 11.1f
C14115 XDAC1.XC64a<0>.XRES4.B AVSS 11.1f
C14116 li_14804_12216# AVSS 0.0299f $ **FLOATING
C14117 li_9184_12216# AVSS 0.0299f $ **FLOATING
C14118 XDAC2.XC64a<0>.XRES1B.B AVSS 8.69f
C14119 XDAC1.XC64a<0>.XRES1B.B AVSS 8.69f
C14120 li_14804_12636# AVSS 0.0299f $ **FLOATING
C14121 XDAC2.XC32a<0>.XRES1A.A AVSS 0.116f
C14122 XDAC1.XC32a<0>.XRES1A.A AVSS 0.116f
C14123 li_9184_12636# AVSS 0.0299f $ **FLOATING
C14124 li_14804_13248# AVSS 0.0311f $ **FLOATING
C14125 li_9184_13248# AVSS 0.0311f $ **FLOATING
C14126 XDAC2.XC32a<0>.XRES16.B AVSS 23.3f
C14127 XDAC1.XC32a<0>.XRES16.B AVSS 23.3f
C14128 li_14804_13860# AVSS 0.031f $ **FLOATING
C14129 li_9184_13860# AVSS 0.031f $ **FLOATING
C14130 XDAC2.XC32a<0>.XRES2.B AVSS 9.11f
C14131 XDAC1.XC32a<0>.XRES2.B AVSS 9.11f
C14132 li_14804_14472# AVSS 0.031f $ **FLOATING
C14133 li_9184_14472# AVSS 0.031f $ **FLOATING
C14134 XDAC2.XC32a<0>.XRES8.B AVSS 15f
C14135 XDAC1.XC32a<0>.XRES8.B AVSS 15f
C14136 li_14804_15084# AVSS 0.0311f $ **FLOATING
C14137 li_9184_15084# AVSS 0.0311f $ **FLOATING
C14138 XDAC2.XC32a<0>.XRES4.B AVSS 11.1f
C14139 XDAC1.XC32a<0>.XRES4.B AVSS 11.1f
C14140 li_14804_15696# AVSS 0.0299f $ **FLOATING
C14141 li_9184_15696# AVSS 0.0299f $ **FLOATING
C14142 XDAC2.XC32a<0>.XRES1B.B AVSS 8.08f
C14143 XDAC1.XC32a<0>.XRES1B.B AVSS 8.08f
C14144 li_14804_16116# AVSS 0.0299f $ **FLOATING
C14145 li_9184_16116# AVSS 0.0299f $ **FLOATING
C14146 XDAC2.XC128a<1>.XRES1A.B AVSS 8.06f
C14147 XDAC1.XC128a<1>.XRES1A.B AVSS 8.06f
C14148 li_14804_16728# AVSS 0.0311f $ **FLOATING
C14149 li_9184_16728# AVSS 0.0311f $ **FLOATING
C14150 XDAC2.XC128a<1>.XRES16.B AVSS 22.8f
C14151 XDAC1.XC128a<1>.XRES16.B AVSS 22.8f
C14152 li_14804_17340# AVSS 0.031f $ **FLOATING
C14153 li_9184_17340# AVSS 0.031f $ **FLOATING
C14154 XDAC2.XC128a<1>.XRES2.B AVSS 9.09f
C14155 XDAC1.XC128a<1>.XRES2.B AVSS 9.09f
C14156 li_14804_17952# AVSS 0.031f $ **FLOATING
C14157 li_9184_17952# AVSS 0.031f $ **FLOATING
C14158 XDAC2.XC128a<1>.XRES8.B AVSS 15f
C14159 XDAC1.XC128a<1>.XRES8.B AVSS 15f
C14160 li_14804_18564# AVSS 0.0311f $ **FLOATING
C14161 li_9184_18564# AVSS 0.0311f $ **FLOATING
C14162 XDAC2.XC128a<1>.XRES4.B AVSS 11.1f
C14163 XDAC1.XC128a<1>.XRES4.B AVSS 11.1f
C14164 li_14804_19176# AVSS 0.0299f $ **FLOATING
C14165 li_9184_19176# AVSS 0.0299f $ **FLOATING
C14166 XDAC2.XC128a<1>.XRES1B.B AVSS 8.07f
C14167 XDAC1.XC128a<1>.XRES1B.B AVSS 8.07f
C14168 li_14804_19596# AVSS 0.0299f $ **FLOATING
C14169 li_9184_19596# AVSS 0.0299f $ **FLOATING
C14170 XDAC2.XC128b<2>.XRES1A.B AVSS 8.06f
C14171 XDAC1.XC128b<2>.XRES1A.B AVSS 8.06f
C14172 li_14804_20208# AVSS 0.0311f $ **FLOATING
C14173 li_9184_20208# AVSS 0.0311f $ **FLOATING
C14174 XDAC2.XC128b<2>.XRES16.B AVSS 22.8f
C14175 XDAC1.XC128b<2>.XRES16.B AVSS 22.8f
C14176 li_14804_20820# AVSS 0.031f $ **FLOATING
C14177 li_9184_20820# AVSS 0.031f $ **FLOATING
C14178 XDAC2.XC128b<2>.XRES2.B AVSS 9.09f
C14179 XDAC1.XC128b<2>.XRES2.B AVSS 9.09f
C14180 li_14804_21432# AVSS 0.031f $ **FLOATING
C14181 li_9184_21432# AVSS 0.031f $ **FLOATING
C14182 XDAC2.XC128b<2>.XRES8.B AVSS 15f
C14183 XDAC1.XC128b<2>.XRES8.B AVSS 15f
C14184 li_14804_22044# AVSS 0.0311f $ **FLOATING
C14185 li_9184_22044# AVSS 0.0311f $ **FLOATING
C14186 XDAC2.XC128b<2>.XRES4.B AVSS 11.1f
C14187 XDAC1.XC128b<2>.XRES4.B AVSS 11.1f
C14188 li_14804_22656# AVSS 0.0299f $ **FLOATING
C14189 li_9184_22656# AVSS 0.0299f $ **FLOATING
C14190 XDAC2.XC128b<2>.XRES1B.B AVSS 8.07f
C14191 XDAC1.XC128b<2>.XRES1B.B AVSS 8.07f
C14192 li_14804_23076# AVSS 0.0299f $ **FLOATING
C14193 li_9184_23076# AVSS 0.0299f $ **FLOATING
C14194 XDAC2.X16ab.XRES1A.B AVSS 8.06f
C14195 XDAC1.X16ab.XRES1A.B AVSS 8.06f
C14196 li_14804_23688# AVSS 0.0311f $ **FLOATING
C14197 li_9184_23688# AVSS 0.0311f $ **FLOATING
C14198 XDAC2.X16ab.XRES16.B AVSS 22.8f
C14199 XDAC1.X16ab.XRES16.B AVSS 22.8f
C14200 li_14804_24300# AVSS 0.031f $ **FLOATING
C14201 li_9184_24300# AVSS 0.031f $ **FLOATING
C14202 XDAC2.X16ab.XRES2.B AVSS 9.09f
C14203 XDAC1.X16ab.XRES2.B AVSS 9.09f
C14204 li_14804_24912# AVSS 0.031f $ **FLOATING
C14205 li_9184_24912# AVSS 0.031f $ **FLOATING
C14206 XDAC2.X16ab.XRES8.B AVSS 15f
C14207 XDAC1.X16ab.XRES8.B AVSS 15f
C14208 li_14804_25524# AVSS 0.0311f $ **FLOATING
C14209 li_9184_25524# AVSS 0.0311f $ **FLOATING
C14210 XDAC2.X16ab.XRES4.B AVSS 11.1f
C14211 XDAC1.X16ab.XRES4.B AVSS 11.1f
C14212 li_14804_26136# AVSS 0.0299f $ **FLOATING
C14213 li_9184_26136# AVSS 0.0299f $ **FLOATING
C14214 XDAC2.X16ab.XRES1B.B AVSS 8.07f
C14215 XDAC1.X16ab.XRES1B.B AVSS 8.07f
C14216 li_14804_26556# AVSS 0.0299f $ **FLOATING
C14217 li_9184_26556# AVSS 0.0299f $ **FLOATING
C14218 XDAC2.XC64b<1>.XRES1A.B AVSS 8.06f
C14219 XDAC1.XC64b<1>.XRES1A.B AVSS 8.06f
C14220 li_14804_27168# AVSS 0.0311f $ **FLOATING
C14221 li_9184_27168# AVSS 0.0311f $ **FLOATING
C14222 XDAC2.XC64b<1>.XRES16.B AVSS 22.8f
C14223 XDAC1.XC64b<1>.XRES16.B AVSS 22.8f
C14224 li_14804_27780# AVSS 0.031f $ **FLOATING
C14225 li_9184_27780# AVSS 0.031f $ **FLOATING
C14226 XDAC2.XC64b<1>.XRES2.B AVSS 9.09f
C14227 XDAC1.XC64b<1>.XRES2.B AVSS 9.09f
C14228 li_14804_28392# AVSS 0.031f $ **FLOATING
C14229 li_9184_28392# AVSS 0.031f $ **FLOATING
C14230 XDAC2.XC64b<1>.XRES8.B AVSS 15f
C14231 XDAC1.XC64b<1>.XRES8.B AVSS 15f
C14232 li_14804_29004# AVSS 0.0311f $ **FLOATING
C14233 li_9184_29004# AVSS 0.0311f $ **FLOATING
C14234 XDAC2.XC64b<1>.XRES4.B AVSS 11.1f
C14235 XDAC1.XC64b<1>.XRES4.B AVSS 11.1f
C14236 li_14804_29616# AVSS 0.0299f $ **FLOATING
C14237 li_9184_29616# AVSS 0.0299f $ **FLOATING
C14238 XDAC2.XC64b<1>.XRES1B.B AVSS 8.07f
C14239 XDAC1.XC64b<1>.XRES1B.B AVSS 8.07f
C14240 li_14804_30036# AVSS 0.0299f $ **FLOATING
C14241 li_9184_30036# AVSS 0.0299f $ **FLOATING
C14242 XDAC2.XC0.XRES1A.B AVSS 8.06f
C14243 XDAC1.XC0.XRES1A.B AVSS 8.06f
C14244 li_14804_30648# AVSS 0.0311f $ **FLOATING
C14245 li_9184_30648# AVSS 0.0311f $ **FLOATING
C14246 XDAC2.XC0.XRES16.B AVSS 22.8f
C14247 XDAC1.XC0.XRES16.B AVSS 22.8f
C14248 li_14804_31260# AVSS 0.031f $ **FLOATING
C14249 li_9184_31260# AVSS 0.031f $ **FLOATING
C14250 XDAC2.XC0.XRES2.B AVSS 9.09f
C14251 XDAC1.XC0.XRES2.B AVSS 9.09f
C14252 li_14804_31872# AVSS 0.031f $ **FLOATING
C14253 li_9184_31872# AVSS 0.031f $ **FLOATING
C14254 XDAC2.XC0.XRES8.B AVSS 15f
C14255 XDAC1.XC0.XRES8.B AVSS 15f
C14256 li_14804_32484# AVSS 0.0311f $ **FLOATING
C14257 li_9184_32484# AVSS 0.0311f $ **FLOATING
C14258 XDAC2.XC0.XRES4.B AVSS 11.1f
C14259 XDAC1.XC0.XRES4.B AVSS 11.1f
C14260 li_14804_33096# AVSS 0.035f $ **FLOATING
C14261 li_9184_33096# AVSS 0.035f $ **FLOATING
C14262 XDAC2.XC0.XRES1B.B AVSS 8.75f
C14263 XDAC1.XC0.XRES1B.B AVSS 8.75f
C14264 a_14960_n18# AVSS 0.0952f $ **FLOATING
C14265 a_13808_n18# AVSS 0.539f $ **FLOATING
C14266 a_12368_n18# AVSS 0.428f $ **FLOATING
C14267 a_11000_n18# AVSS 0.427f $ **FLOATING
C14268 a_9560_n18# AVSS 0.54f $ **FLOATING
C14269 a_8408_n18# AVSS 0.0952f $ **FLOATING
C14270 a_14960_334# AVSS 0.00282f $ **FLOATING
C14271 a_13808_334# AVSS 0.488f $ **FLOATING
C14272 a_12368_334# AVSS 0.353f $ **FLOATING
C14273 a_11000_334# AVSS 0.353f $ **FLOATING
C14274 a_9560_334# AVSS 0.487f $ **FLOATING
C14275 a_8408_334# AVSS 0.00282f $ **FLOATING
C14276 CK_SAMPLE_BSSW AVSS 28.3f
C14277 a_14960_686# AVSS 0.00275f $ **FLOATING
C14278 a_13808_686# AVSS 0.365f $ **FLOATING
C14279 a_12368_686# AVSS 0.352f $ **FLOATING
C14280 a_11000_686# AVSS 0.352f $ **FLOATING
C14281 a_9560_686# AVSS 0.365f $ **FLOATING
C14282 a_8408_686# AVSS 0.00275f $ **FLOATING
C14283 a_14960_1038# AVSS 0.00291f $ **FLOATING
C14284 a_13808_1038# AVSS 0.414f $ **FLOATING
C14285 a_12368_1038# AVSS 0.352f $ **FLOATING
C14286 a_11000_1038# AVSS 0.352f $ **FLOATING
C14287 a_9560_1038# AVSS 0.414f $ **FLOATING
C14288 a_8408_1038# AVSS 0.00291f $ **FLOATING
C14289 a_14960_1390# AVSS 0.00269f $ **FLOATING
C14290 a_13808_1390# AVSS 0.363f $ **FLOATING
C14291 a_12368_1390# AVSS 0.354f $ **FLOATING
C14292 a_11000_1390# AVSS 0.354f $ **FLOATING
C14293 a_9560_1390# AVSS 0.363f $ **FLOATING
C14294 a_8408_1390# AVSS 0.00269f $ **FLOATING
C14295 XB2.XA3.MN1.D AVSS 52.2f
C14296 XB2.XA3.MN0.S AVSS 0.813f
C14297 XB1.XA3.MN1.D AVSS 52.2f
C14298 XB1.XA3.MN0.S AVSS 0.813f
C14299 a_14960_1742# AVSS 0.00276f $ **FLOATING
C14300 a_13808_1742# AVSS 0.382f $ **FLOATING
C14301 a_12368_1742# AVSS 0.352f $ **FLOATING
C14302 a_11000_1742# AVSS 0.352f $ **FLOATING
C14303 a_9560_1742# AVSS 0.382f $ **FLOATING
C14304 a_8408_1742# AVSS 0.00276f $ **FLOATING
C14305 XB2.XA0.MP0.D AVSS 2.63f
C14306 XB1.XA0.MP0.D AVSS 2.63f
C14307 a_14960_2094# AVSS 0.00269f $ **FLOATING
C14308 a_13808_2094# AVSS 0.363f $ **FLOATING
C14309 a_12368_2094# AVSS 0.352f $ **FLOATING
C14310 a_11000_2094# AVSS 0.352f $ **FLOATING
C14311 a_9560_2094# AVSS 0.363f $ **FLOATING
C14312 a_8408_2094# AVSS 0.00269f $ **FLOATING
C14313 XB2.XA4.MP0.D AVSS 49f
C14314 XB2.XA4.MN0.D AVSS 0.162f
C14315 XB2.M1.G AVSS 3.18f
C14316 XB1.XA4.MN0.D AVSS 0.162f
C14317 XB1.XA4.MP0.D AVSS 49f
C14318 XB1.M1.G AVSS 3.12f
C14319 a_14960_2446# AVSS 0.00276f $ **FLOATING
C14320 a_13808_2446# AVSS 0.382f $ **FLOATING
C14321 a_12368_2446# AVSS 0.352f $ **FLOATING
C14322 a_11000_2446# AVSS 0.352f $ **FLOATING
C14323 a_9560_2446# AVSS 0.382f $ **FLOATING
C14324 a_8408_2446# AVSS 0.00276f $ **FLOATING
C14325 XB2.XA1.MP0.D AVSS 0.941f
C14326 SAR_IN AVSS 1.81f
C14327 XB2.XA1.MN0.D AVSS 0.786f
C14328 SAR_IP AVSS 1.81f
C14329 XB1.XA1.MN0.D AVSS 0.786f
C14330 XB1.XA1.MP0.D AVSS 0.941f
C14331 a_14960_2798# AVSS 0.00276f $ **FLOATING
C14332 a_13808_2798# AVSS 0.467f $ **FLOATING
C14333 a_12368_2798# AVSS 0.423f $ **FLOATING
C14334 a_11000_2798# AVSS 0.424f $ **FLOATING
C14335 a_9560_2798# AVSS 0.468f $ **FLOATING
C14336 a_8408_2798# AVSS 0.00276f $ **FLOATING
C14337 a_14960_3150# AVSS 0.00276f $ **FLOATING
C14338 a_13808_3150# AVSS 0.49f $ **FLOATING
C14339 XB2.XA2.MN0.G AVSS 0.591f
C14340 a_14960_3502# AVSS 0.00276f $ **FLOATING
C14341 a_13808_3502# AVSS 0.468f $ **FLOATING
C14342 a_14960_3854# AVSS 0.0907f $ **FLOATING
C14343 a_13808_3854# AVSS 0.538f $ **FLOATING
C14344 a_9560_3150# AVSS 0.489f $ **FLOATING
C14345 a_8408_3150# AVSS 0.00276f $ **FLOATING
C14346 XB1.XA2.MN0.G AVSS 0.591f
C14347 a_9560_3502# AVSS 0.47f $ **FLOATING
C14348 a_8408_3502# AVSS 0.00276f $ **FLOATING
C14349 a_9560_3854# AVSS 0.537f $ **FLOATING
C14350 a_8408_3854# AVSS 0.0907f $ **FLOATING
C14351 a_23600_39876# AVSS 0.529f $ **FLOATING
C14352 a_22448_39876# AVSS 0.0889f $ **FLOATING
C14353 a_21080_39876# AVSS 0.0889f $ **FLOATING
C14354 a_19928_39876# AVSS 0.528f $ **FLOATING
C14355 a_18560_39876# AVSS 0.529f $ **FLOATING
C14356 a_17408_39876# AVSS 0.0888f $ **FLOATING
C14357 a_16040_39876# AVSS 0.0888f $ **FLOATING
C14358 a_14888_39876# AVSS 0.528f $ **FLOATING
C14359 a_13520_39876# AVSS 0.529f $ **FLOATING
C14360 a_12368_39876# AVSS 0.0888f $ **FLOATING
C14361 a_11000_39876# AVSS 0.0888f $ **FLOATING
C14362 a_9848_39876# AVSS 0.527f $ **FLOATING
C14363 a_8480_39876# AVSS 0.528f $ **FLOATING
C14364 a_7328_39876# AVSS 0.0888f $ **FLOATING
C14365 a_5960_39876# AVSS 0.0888f $ **FLOATING
C14366 a_4808_39876# AVSS 0.527f $ **FLOATING
C14367 a_3440_39876# AVSS 0.528f $ **FLOATING
C14368 a_2288_39876# AVSS 0.0888f $ **FLOATING
C14369 a_920_39876# AVSS 0.0888f $ **FLOATING
C14370 a_n232_39876# AVSS 0.528f $ **FLOATING
C14371 a_23600_40228# AVSS 0.487f $ **FLOATING
C14372 a_22448_40228# AVSS 0.00159f $ **FLOATING
C14373 a_21080_40228# AVSS 0.00159f $ **FLOATING
C14374 a_19928_40228# AVSS 0.469f $ **FLOATING
C14375 a_18560_40228# AVSS 0.463f $ **FLOATING
C14376 a_17408_40228# AVSS 0.00131f $ **FLOATING
C14377 a_16040_40228# AVSS 0.00131f $ **FLOATING
C14378 a_14888_40228# AVSS 0.469f $ **FLOATING
C14379 a_13520_40228# AVSS 0.463f $ **FLOATING
C14380 a_12368_40228# AVSS 0.00131f $ **FLOATING
C14381 a_11000_40228# AVSS 0.00131f $ **FLOATING
C14382 a_9848_40228# AVSS 0.468f $ **FLOATING
C14383 a_8480_40228# AVSS 0.461f $ **FLOATING
C14384 a_7328_40228# AVSS 0.00131f $ **FLOATING
C14385 a_5960_40228# AVSS 0.00131f $ **FLOATING
C14386 a_4808_40228# AVSS 0.468f $ **FLOATING
C14387 a_3440_40228# AVSS 0.461f $ **FLOATING
C14388 a_2288_40228# AVSS 0.00131f $ **FLOATING
C14389 a_920_40228# AVSS 0.00131f $ **FLOATING
C14390 a_n232_40228# AVSS 0.469f $ **FLOATING
C14391 a_23600_40580# AVSS 0.363f $ **FLOATING
C14392 a_22448_40580# AVSS 0.00152f $ **FLOATING
C14393 a_21080_40580# AVSS 0.00152f $ **FLOATING
C14394 a_19928_40580# AVSS 0.385f $ **FLOATING
C14395 a_18560_40580# AVSS 0.384f $ **FLOATING
C14396 a_17408_40580# AVSS 0.00125f $ **FLOATING
C14397 a_16040_40580# AVSS 0.00125f $ **FLOATING
C14398 a_14888_40580# AVSS 0.385f $ **FLOATING
C14399 a_13520_40580# AVSS 0.384f $ **FLOATING
C14400 a_12368_40580# AVSS 0.00125f $ **FLOATING
C14401 a_11000_40580# AVSS 0.00125f $ **FLOATING
C14402 a_9848_40580# AVSS 0.385f $ **FLOATING
C14403 a_8480_40580# AVSS 0.382f $ **FLOATING
C14404 a_7328_40580# AVSS 0.00125f $ **FLOATING
C14405 a_5960_40580# AVSS 0.00125f $ **FLOATING
C14406 a_4808_40580# AVSS 0.384f $ **FLOATING
C14407 a_3440_40580# AVSS 0.382f $ **FLOATING
C14408 a_2288_40580# AVSS 0.00125f $ **FLOATING
C14409 a_920_40580# AVSS 0.00125f $ **FLOATING
C14410 a_n232_40580# AVSS 0.385f $ **FLOATING
C14411 a_23600_40932# AVSS 0.358f $ **FLOATING
C14412 a_22448_40932# AVSS 0.00152f $ **FLOATING
C14413 a_21080_40932# AVSS 0.00148f $ **FLOATING
C14414 a_19928_40932# AVSS 0.369f $ **FLOATING
C14415 a_18560_40932# AVSS 0.367f $ **FLOATING
C14416 a_17408_40932# AVSS 0.00125f $ **FLOATING
C14417 a_16040_40932# AVSS 0.00125f $ **FLOATING
C14418 a_14888_40932# AVSS 0.369f $ **FLOATING
C14419 a_13520_40932# AVSS 0.367f $ **FLOATING
C14420 a_12368_40932# AVSS 0.00125f $ **FLOATING
C14421 a_11000_40932# AVSS 0.00125f $ **FLOATING
C14422 a_9848_40932# AVSS 0.368f $ **FLOATING
C14423 a_8480_40932# AVSS 0.366f $ **FLOATING
C14424 a_7328_40932# AVSS 0.00125f $ **FLOATING
C14425 a_5960_40932# AVSS 0.00125f $ **FLOATING
C14426 a_4808_40932# AVSS 0.368f $ **FLOATING
C14427 a_3440_40932# AVSS 0.366f $ **FLOATING
C14428 a_2288_40932# AVSS 0.00125f $ **FLOATING
C14429 a_920_40932# AVSS 0.00125f $ **FLOATING
C14430 a_n232_40932# AVSS 0.369f $ **FLOATING
C14431 XA8.XA1.XA1.MN0.D AVSS 0.478f
C14432 XA7.XA1.XA1.MN0.D AVSS 0.451f
C14433 XA6.XA1.XA1.MN0.D AVSS 0.474f
C14434 XA5.XA1.XA1.MN0.D AVSS 0.451f
C14435 XA4.XA1.XA1.MN0.D AVSS 0.474f
C14436 XA3.XA1.XA1.MN0.D AVSS 0.451f
C14437 XA2.XA1.XA1.MN0.D AVSS 0.474f
C14438 XA1.XA1.XA1.MN0.D AVSS 0.451f
C14439 XA0.XA1.XA1.MN0.D AVSS 0.474f
C14440 a_23600_41284# AVSS 0.357f $ **FLOATING
C14441 a_22448_41284# AVSS 0.00152f $ **FLOATING
C14442 a_21080_41284# AVSS 0.00148f $ **FLOATING
C14443 a_19928_41284# AVSS 0.404f $ **FLOATING
C14444 a_18560_41284# AVSS 0.404f $ **FLOATING
C14445 a_17408_41284# AVSS 0.00125f $ **FLOATING
C14446 a_16040_41284# AVSS 0.00125f $ **FLOATING
C14447 a_14888_41284# AVSS 0.404f $ **FLOATING
C14448 a_13520_41284# AVSS 0.404f $ **FLOATING
C14449 a_12368_41284# AVSS 0.00125f $ **FLOATING
C14450 a_11000_41284# AVSS 0.00125f $ **FLOATING
C14451 a_9848_41284# AVSS 0.403f $ **FLOATING
C14452 a_8480_41284# AVSS 0.402f $ **FLOATING
C14453 a_7328_41284# AVSS 0.00125f $ **FLOATING
C14454 a_5960_41284# AVSS 0.00125f $ **FLOATING
C14455 a_4808_41284# AVSS 0.403f $ **FLOATING
C14456 a_3440_41284# AVSS 0.402f $ **FLOATING
C14457 a_2288_41284# AVSS 0.00125f $ **FLOATING
C14458 a_920_41284# AVSS 0.00125f $ **FLOATING
C14459 a_n232_41284# AVSS 0.404f $ **FLOATING
C14460 XA8.XA1.XA1.MP2.D AVSS 0.00324f
C14461 XA8.XA1.XA1.MN0.S AVSS 0.745f
C14462 XA7.XA1.XA1.MP2.D AVSS 0.00324f
C14463 XA7.XA1.XA1.MN0.S AVSS 0.728f
C14464 XA6.XA1.XA1.MP2.D AVSS 0.00324f
C14465 XA6.XA1.XA1.MN0.S AVSS 0.738f
C14466 XA5.XA1.XA1.MP2.D AVSS 0.00324f
C14467 XA5.XA1.XA1.MN0.S AVSS 0.728f
C14468 XA4.XA1.XA1.MP2.D AVSS 0.00324f
C14469 XA4.XA1.XA1.MN0.S AVSS 0.737f
C14470 XA3.XA1.XA1.MP2.D AVSS 0.00324f
C14471 XA3.XA1.XA1.MN0.S AVSS 0.725f
C14472 XA2.XA1.XA1.MP2.D AVSS 0.00324f
C14473 XA2.XA1.XA1.MN0.S AVSS 0.736f
C14474 XA1.XA1.XA1.MP2.D AVSS 0.00324f
C14475 XA1.XA1.XA1.MN0.S AVSS 0.724f
C14476 XA0.XA1.XA1.MP2.D AVSS 0.00324f
C14477 XA0.XA1.XA1.MN0.S AVSS 0.738f
C14478 a_23600_41636# AVSS 0.357f $ **FLOATING
C14479 a_22448_41636# AVSS 0.00152f $ **FLOATING
C14480 a_21080_41636# AVSS 0.00152f $ **FLOATING
C14481 a_19928_41636# AVSS 0.386f $ **FLOATING
C14482 a_18560_41636# AVSS 0.386f $ **FLOATING
C14483 a_17408_41636# AVSS 0.00125f $ **FLOATING
C14484 a_16040_41636# AVSS 0.00125f $ **FLOATING
C14485 a_14888_41636# AVSS 0.386f $ **FLOATING
C14486 a_13520_41636# AVSS 0.386f $ **FLOATING
C14487 a_12368_41636# AVSS 0.00125f $ **FLOATING
C14488 a_11000_41636# AVSS 0.00125f $ **FLOATING
C14489 a_9848_41636# AVSS 0.385f $ **FLOATING
C14490 a_8480_41636# AVSS 0.384f $ **FLOATING
C14491 a_7328_41636# AVSS 0.00125f $ **FLOATING
C14492 a_5960_41636# AVSS 0.00125f $ **FLOATING
C14493 a_4808_41636# AVSS 0.385f $ **FLOATING
C14494 a_3440_41636# AVSS 0.384f $ **FLOATING
C14495 a_2288_41636# AVSS 0.00125f $ **FLOATING
C14496 a_920_41636# AVSS 0.00125f $ **FLOATING
C14497 a_n232_41636# AVSS 0.386f $ **FLOATING
C14498 a_23600_41988# AVSS 0.357f $ **FLOATING
C14499 a_22448_41988# AVSS 0.00152f $ **FLOATING
C14500 a_21080_41988# AVSS 0.00152f $ **FLOATING
C14501 a_19928_41988# AVSS 0.385f $ **FLOATING
C14502 a_18560_41988# AVSS 0.386f $ **FLOATING
C14503 a_17408_41988# AVSS 0.00125f $ **FLOATING
C14504 a_16040_41988# AVSS 0.00125f $ **FLOATING
C14505 a_14888_41988# AVSS 0.386f $ **FLOATING
C14506 a_13520_41988# AVSS 0.386f $ **FLOATING
C14507 a_12368_41988# AVSS 0.00125f $ **FLOATING
C14508 a_11000_41988# AVSS 0.00125f $ **FLOATING
C14509 a_9848_41988# AVSS 0.385f $ **FLOATING
C14510 a_8480_41988# AVSS 0.384f $ **FLOATING
C14511 a_7328_41988# AVSS 0.00125f $ **FLOATING
C14512 a_5960_41988# AVSS 0.00125f $ **FLOATING
C14513 a_4808_41988# AVSS 0.385f $ **FLOATING
C14514 a_3440_41988# AVSS 0.384f $ **FLOATING
C14515 a_2288_41988# AVSS 0.00125f $ **FLOATING
C14516 a_920_41988# AVSS 0.00125f $ **FLOATING
C14517 a_n232_41988# AVSS 0.386f $ **FLOATING
C14518 a_23600_42340# AVSS 0.36f $ **FLOATING
C14519 a_22448_42340# AVSS 0.00152f $ **FLOATING
C14520 a_21080_42340# AVSS 0.00152f $ **FLOATING
C14521 a_19928_42340# AVSS 0.36f $ **FLOATING
C14522 a_18560_42340# AVSS 0.36f $ **FLOATING
C14523 a_17408_42340# AVSS 0.00125f $ **FLOATING
C14524 a_16040_42340# AVSS 0.00125f $ **FLOATING
C14525 a_14888_42340# AVSS 0.361f $ **FLOATING
C14526 a_13520_42340# AVSS 0.36f $ **FLOATING
C14527 a_12368_42340# AVSS 0.00125f $ **FLOATING
C14528 a_11000_42340# AVSS 0.00125f $ **FLOATING
C14529 a_9848_42340# AVSS 0.36f $ **FLOATING
C14530 a_8480_42340# AVSS 0.359f $ **FLOATING
C14531 a_7328_42340# AVSS 0.00125f $ **FLOATING
C14532 a_5960_42340# AVSS 0.00125f $ **FLOATING
C14533 a_4808_42340# AVSS 0.36f $ **FLOATING
C14534 a_3440_42340# AVSS 0.359f $ **FLOATING
C14535 a_2288_42340# AVSS 0.00125f $ **FLOATING
C14536 a_920_42340# AVSS 0.00125f $ **FLOATING
C14537 a_n232_42340# AVSS 0.361f $ **FLOATING
C14538 XA20.XA1.MN0.D AVSS 0.946f
C14539 XA8.XA1.XA4.MP0.D AVSS 0.00883f
C14540 XA8.XA1.XA4.MN0.D AVSS 0.134f
C14541 XA7.XA1.XA4.MN0.D AVSS 0.139f
C14542 XA7.XA1.XA4.MP0.D AVSS 0.00883f
C14543 XA6.XA1.XA4.MP0.D AVSS 0.00883f
C14544 XA6.XA1.XA4.MN0.D AVSS 0.139f
C14545 XA5.XA1.XA4.MN0.D AVSS 0.139f
C14546 XA5.XA1.XA4.MP0.D AVSS 0.00883f
C14547 XA4.XA1.XA4.MP0.D AVSS 0.00883f
C14548 XA4.XA1.XA4.MN0.D AVSS 0.139f
C14549 XA3.XA1.XA4.MN0.D AVSS 0.139f
C14550 XA3.XA1.XA4.MP0.D AVSS 0.00883f
C14551 XA2.XA1.XA4.MP0.D AVSS 0.00883f
C14552 XA2.XA1.XA4.MN0.D AVSS 0.139f
C14553 XA1.XA1.XA4.MN0.D AVSS 0.139f
C14554 XA1.XA1.XA4.MP0.D AVSS 0.00883f
C14555 XA0.XA1.XA4.MP0.D AVSS 0.00883f
C14556 XA0.XA1.XA4.MN0.D AVSS 0.139f
C14557 a_23600_42692# AVSS 0.381f $ **FLOATING
C14558 a_22448_42692# AVSS 0.00152f $ **FLOATING
C14559 a_21080_42692# AVSS 0.00152f $ **FLOATING
C14560 a_19928_42692# AVSS 0.358f $ **FLOATING
C14561 a_18560_42692# AVSS 0.357f $ **FLOATING
C14562 a_17408_42692# AVSS 0.00125f $ **FLOATING
C14563 a_16040_42692# AVSS 0.00125f $ **FLOATING
C14564 a_14888_42692# AVSS 0.357f $ **FLOATING
C14565 a_13520_42692# AVSS 0.357f $ **FLOATING
C14566 a_12368_42692# AVSS 0.00125f $ **FLOATING
C14567 a_11000_42692# AVSS 0.00125f $ **FLOATING
C14568 a_9848_42692# AVSS 0.356f $ **FLOATING
C14569 a_8480_42692# AVSS 0.355f $ **FLOATING
C14570 a_7328_42692# AVSS 0.00125f $ **FLOATING
C14571 a_5960_42692# AVSS 0.00125f $ **FLOATING
C14572 a_4808_42692# AVSS 0.356f $ **FLOATING
C14573 a_3440_42692# AVSS 0.355f $ **FLOATING
C14574 a_2288_42692# AVSS 0.00125f $ **FLOATING
C14575 a_920_42692# AVSS 0.00125f $ **FLOATING
C14576 a_n232_42692# AVSS 0.357f $ **FLOATING
C14577 XA8.XA1.XA4.MP1.D AVSS 0.00883f
C14578 XA8.XA1.XA4.MN1.D AVSS 0.0813f
C14579 XA7.XA1.XA4.MN1.D AVSS 0.0736f
C14580 XA7.XA1.XA4.MP1.D AVSS 0.00883f
C14581 XA6.XA1.XA4.MP1.D AVSS 0.00883f
C14582 XA6.XA1.XA4.MN1.D AVSS 0.0736f
C14583 XA5.XA1.XA4.MN1.D AVSS 0.0736f
C14584 XA5.XA1.XA4.MP1.D AVSS 0.00883f
C14585 XA4.XA1.XA4.MP1.D AVSS 0.00883f
C14586 XA4.XA1.XA4.MN1.D AVSS 0.0736f
C14587 XA3.XA1.XA4.MN1.D AVSS 0.0736f
C14588 XA3.XA1.XA4.MP1.D AVSS 0.00883f
C14589 XA2.XA1.XA4.MP1.D AVSS 0.00883f
C14590 XA2.XA1.XA4.MN1.D AVSS 0.0736f
C14591 XA1.XA1.XA4.MN1.D AVSS 0.0736f
C14592 XA1.XA1.XA4.MP1.D AVSS 0.00883f
C14593 XA0.XA1.XA4.MP1.D AVSS 0.00883f
C14594 XA0.XA1.XA4.MN1.D AVSS 0.0736f
C14595 a_23600_43044# AVSS 0.361f $ **FLOATING
C14596 a_22448_43044# AVSS 0.00152f $ **FLOATING
C14597 a_21080_43044# AVSS 0.00152f $ **FLOATING
C14598 a_19928_43044# AVSS 0.38f $ **FLOATING
C14599 a_18560_43044# AVSS 0.38f $ **FLOATING
C14600 a_17408_43044# AVSS 0.00125f $ **FLOATING
C14601 a_16040_43044# AVSS 0.00125f $ **FLOATING
C14602 a_14888_43044# AVSS 0.38f $ **FLOATING
C14603 a_13520_43044# AVSS 0.38f $ **FLOATING
C14604 a_12368_43044# AVSS 0.00125f $ **FLOATING
C14605 a_11000_43044# AVSS 0.00125f $ **FLOATING
C14606 a_9848_43044# AVSS 0.379f $ **FLOATING
C14607 a_8480_43044# AVSS 0.378f $ **FLOATING
C14608 a_7328_43044# AVSS 0.00125f $ **FLOATING
C14609 a_5960_43044# AVSS 0.00125f $ **FLOATING
C14610 a_4808_43044# AVSS 0.379f $ **FLOATING
C14611 a_3440_43044# AVSS 0.378f $ **FLOATING
C14612 a_2288_43044# AVSS 0.00125f $ **FLOATING
C14613 a_920_43044# AVSS 0.00125f $ **FLOATING
C14614 a_n232_43044# AVSS 0.38f $ **FLOATING
C14615 a_23600_43396# AVSS 0.358f $ **FLOATING
C14616 a_22448_43396# AVSS 0.00152f $ **FLOATING
C14617 a_21080_43396# AVSS 0.00152f $ **FLOATING
C14618 a_19928_43396# AVSS 0.362f $ **FLOATING
C14619 a_18560_43396# AVSS 0.363f $ **FLOATING
C14620 a_17408_43396# AVSS 0.00125f $ **FLOATING
C14621 a_16040_43396# AVSS 0.00125f $ **FLOATING
C14622 a_14888_43396# AVSS 0.363f $ **FLOATING
C14623 a_13520_43396# AVSS 0.363f $ **FLOATING
C14624 a_12368_43396# AVSS 0.00125f $ **FLOATING
C14625 a_11000_43396# AVSS 0.00125f $ **FLOATING
C14626 a_9848_43396# AVSS 0.362f $ **FLOATING
C14627 a_8480_43396# AVSS 0.361f $ **FLOATING
C14628 a_7328_43396# AVSS 0.00125f $ **FLOATING
C14629 a_5960_43396# AVSS 0.00125f $ **FLOATING
C14630 a_4808_43396# AVSS 0.362f $ **FLOATING
C14631 a_3440_43396# AVSS 0.361f $ **FLOATING
C14632 a_2288_43396# AVSS 0.00125f $ **FLOATING
C14633 a_920_43396# AVSS 0.00125f $ **FLOATING
C14634 a_n232_43396# AVSS 0.363f $ **FLOATING
C14635 XA8.XA1.XA5.MP0.D AVSS 0.00882f
C14636 XA8.XA1.XA5.MN0.D AVSS 0.134f
C14637 XA8.XA1.XA2.MP0.D AVSS 1.42f
C14638 XA7.XA1.XA5.MN0.D AVSS 0.15f
C14639 XA7.XA1.XA5.MP0.D AVSS 0.00883f
C14640 XA7.XA1.XA2.MP0.D AVSS 1.41f
C14641 XA6.XA1.XA5.MP0.D AVSS 0.00883f
C14642 XA6.XA1.XA5.MN0.D AVSS 0.15f
C14643 XA6.XA1.XA2.MP0.D AVSS 1.41f
C14644 XA5.XA1.XA5.MN0.D AVSS 0.15f
C14645 XA5.XA1.XA5.MP0.D AVSS 0.00883f
C14646 XA5.XA1.XA2.MP0.D AVSS 1.41f
C14647 XA4.XA1.XA5.MP0.D AVSS 0.00883f
C14648 XA4.XA1.XA5.MN0.D AVSS 0.15f
C14649 XA4.XA1.XA2.MP0.D AVSS 1.41f
C14650 XA3.XA1.XA5.MN0.D AVSS 0.15f
C14651 XA3.XA1.XA5.MP0.D AVSS 0.00883f
C14652 XA3.XA1.XA2.MP0.D AVSS 1.41f
C14653 XA2.XA1.XA5.MP0.D AVSS 0.00883f
C14654 XA2.XA1.XA5.MN0.D AVSS 0.15f
C14655 XA2.XA1.XA2.MP0.D AVSS 1.41f
C14656 XA1.XA1.XA5.MN0.D AVSS 0.15f
C14657 XA1.XA1.XA5.MP0.D AVSS 0.00883f
C14658 XA1.XA1.XA2.MP0.D AVSS 1.4f
C14659 XA0.XA1.XA5.MP0.D AVSS 0.00883f
C14660 XA0.XA1.XA5.MN0.D AVSS 0.15f
C14661 XA0.XA1.XA2.MP0.D AVSS 1.41f
C14662 a_23600_43748# AVSS 0.357f $ **FLOATING
C14663 a_22448_43748# AVSS 0.00152f $ **FLOATING
C14664 a_21080_43748# AVSS 0.00152f $ **FLOATING
C14665 a_19928_43748# AVSS 0.359f $ **FLOATING
C14666 a_18560_43748# AVSS 0.36f $ **FLOATING
C14667 a_17408_43748# AVSS 0.00125f $ **FLOATING
C14668 a_16040_43748# AVSS 0.00125f $ **FLOATING
C14669 a_14888_43748# AVSS 0.36f $ **FLOATING
C14670 a_13520_43748# AVSS 0.36f $ **FLOATING
C14671 a_12368_43748# AVSS 0.00125f $ **FLOATING
C14672 a_11000_43748# AVSS 0.00125f $ **FLOATING
C14673 a_9848_43748# AVSS 0.359f $ **FLOATING
C14674 a_8480_43748# AVSS 0.359f $ **FLOATING
C14675 a_7328_43748# AVSS 0.00125f $ **FLOATING
C14676 a_5960_43748# AVSS 0.00125f $ **FLOATING
C14677 a_4808_43748# AVSS 0.359f $ **FLOATING
C14678 a_3440_43748# AVSS 0.358f $ **FLOATING
C14679 a_2288_43748# AVSS 0.00125f $ **FLOATING
C14680 a_920_43748# AVSS 0.00125f $ **FLOATING
C14681 a_n232_43748# AVSS 0.36f $ **FLOATING
C14682 XA8.XA1.XA5.MP1.D AVSS 0.00893f
C14683 XA8.XA1.XA5.MN1.D AVSS 0.108f
C14684 XA7.XA1.XA5.MN1.D AVSS 0.113f
C14685 XA7.XA1.XA5.MP1.D AVSS 0.00893f
C14686 XA6.XA1.XA5.MP1.D AVSS 0.00893f
C14687 XA6.XA1.XA5.MN1.D AVSS 0.113f
C14688 XA5.XA1.XA5.MN1.D AVSS 0.113f
C14689 XA5.XA1.XA5.MP1.D AVSS 0.00893f
C14690 XA4.XA1.XA5.MP1.D AVSS 0.00893f
C14691 XA4.XA1.XA5.MN1.D AVSS 0.113f
C14692 XA3.XA1.XA5.MN1.D AVSS 0.113f
C14693 XA3.XA1.XA5.MP1.D AVSS 0.00893f
C14694 XA2.XA1.XA5.MP1.D AVSS 0.00893f
C14695 XA2.XA1.XA5.MN1.D AVSS 0.113f
C14696 XA1.XA1.XA5.MN1.D AVSS 0.113f
C14697 XA1.XA1.XA5.MP1.D AVSS 0.00893f
C14698 XA0.XA1.XA5.MP1.D AVSS 0.00893f
C14699 XA0.XA1.XA5.MN1.D AVSS 0.113f
C14700 EN AVSS 8.08f
C14701 a_23600_44100# AVSS 0.357f $ **FLOATING
C14702 a_22448_44100# AVSS 0.00148f $ **FLOATING
C14703 a_21080_44100# AVSS 0.00159f $ **FLOATING
C14704 a_19928_44100# AVSS 0.382f $ **FLOATING
C14705 a_18560_44100# AVSS 0.382f $ **FLOATING
C14706 a_17408_44100# AVSS 0.00131f $ **FLOATING
C14707 a_16040_44100# AVSS 0.00131f $ **FLOATING
C14708 a_14888_44100# AVSS 0.382f $ **FLOATING
C14709 a_13520_44100# AVSS 0.382f $ **FLOATING
C14710 a_12368_44100# AVSS 0.00131f $ **FLOATING
C14711 a_11000_44100# AVSS 0.00131f $ **FLOATING
C14712 a_9848_44100# AVSS 0.382f $ **FLOATING
C14713 a_8480_44100# AVSS 0.381f $ **FLOATING
C14714 a_7328_44100# AVSS 0.00131f $ **FLOATING
C14715 a_5960_44100# AVSS 0.00131f $ **FLOATING
C14716 a_4808_44100# AVSS 0.381f $ **FLOATING
C14717 a_3440_44100# AVSS 0.38f $ **FLOATING
C14718 a_2288_44100# AVSS 0.00131f $ **FLOATING
C14719 a_920_44100# AVSS 0.00131f $ **FLOATING
C14720 a_n232_44100# AVSS 0.382f $ **FLOATING
C14721 a_23600_44452# AVSS 0.357f $ **FLOATING
C14722 a_22448_44452# AVSS 0.00148f $ **FLOATING
C14723 a_21080_44452# AVSS 0.00152f $ **FLOATING
C14724 a_19928_44452# AVSS 0.366f $ **FLOATING
C14725 a_18560_44452# AVSS 0.366f $ **FLOATING
C14726 a_17408_44452# AVSS 0.00125f $ **FLOATING
C14727 a_16040_44452# AVSS 0.00125f $ **FLOATING
C14728 a_14888_44452# AVSS 0.366f $ **FLOATING
C14729 a_13520_44452# AVSS 0.366f $ **FLOATING
C14730 a_12368_44452# AVSS 0.00125f $ **FLOATING
C14731 a_11000_44452# AVSS 0.00125f $ **FLOATING
C14732 a_9848_44452# AVSS 0.365f $ **FLOATING
C14733 a_8480_44452# AVSS 0.364f $ **FLOATING
C14734 a_7328_44452# AVSS 0.00125f $ **FLOATING
C14735 a_5960_44452# AVSS 0.00125f $ **FLOATING
C14736 a_4808_44452# AVSS 0.365f $ **FLOATING
C14737 a_3440_44452# AVSS 0.364f $ **FLOATING
C14738 a_2288_44452# AVSS 0.00125f $ **FLOATING
C14739 a_920_44452# AVSS 0.00125f $ **FLOATING
C14740 a_n232_44452# AVSS 0.366f $ **FLOATING
C14741 SARP AVSS 0.305p
C14742 a_23600_44804# AVSS 0.359f $ **FLOATING
C14743 a_22448_44804# AVSS 0.00148f $ **FLOATING
C14744 a_21080_44804# AVSS 0.00152f $ **FLOATING
C14745 a_19928_44804# AVSS 0.414f $ **FLOATING
C14746 a_18560_44804# AVSS 0.414f $ **FLOATING
C14747 a_17408_44804# AVSS 0.00125f $ **FLOATING
C14748 a_16040_44804# AVSS 0.00125f $ **FLOATING
C14749 a_14888_44804# AVSS 0.414f $ **FLOATING
C14750 a_13520_44804# AVSS 0.414f $ **FLOATING
C14751 a_12368_44804# AVSS 0.00125f $ **FLOATING
C14752 a_11000_44804# AVSS 0.00125f $ **FLOATING
C14753 a_9848_44804# AVSS 0.413f $ **FLOATING
C14754 a_8480_44804# AVSS 0.413f $ **FLOATING
C14755 a_7328_44804# AVSS 0.00125f $ **FLOATING
C14756 a_5960_44804# AVSS 0.00125f $ **FLOATING
C14757 a_4808_44804# AVSS 0.413f $ **FLOATING
C14758 a_3440_44804# AVSS 0.412f $ **FLOATING
C14759 a_2288_44804# AVSS 0.00125f $ **FLOATING
C14760 a_920_44804# AVSS 0.00125f $ **FLOATING
C14761 a_n232_44804# AVSS 0.414f $ **FLOATING
C14762 XA20.XA2.MN1.D AVSS 0.573f
C14763 a_23600_45156# AVSS 0.38f $ **FLOATING
C14764 a_22448_45156# AVSS 0.00152f $ **FLOATING
C14765 a_21080_45156# AVSS 0.00152f $ **FLOATING
C14766 a_19928_45156# AVSS 0.366f $ **FLOATING
C14767 a_18560_45156# AVSS 0.366f $ **FLOATING
C14768 a_17408_45156# AVSS 0.00125f $ **FLOATING
C14769 a_16040_45156# AVSS 0.00125f $ **FLOATING
C14770 a_14888_45156# AVSS 0.366f $ **FLOATING
C14771 a_13520_45156# AVSS 0.366f $ **FLOATING
C14772 a_12368_45156# AVSS 0.00125f $ **FLOATING
C14773 a_11000_45156# AVSS 0.00125f $ **FLOATING
C14774 a_9848_45156# AVSS 0.365f $ **FLOATING
C14775 a_8480_45156# AVSS 0.364f $ **FLOATING
C14776 a_7328_45156# AVSS 0.00125f $ **FLOATING
C14777 a_5960_45156# AVSS 0.00125f $ **FLOATING
C14778 a_4808_45156# AVSS 0.365f $ **FLOATING
C14779 a_3440_45156# AVSS 0.364f $ **FLOATING
C14780 a_2288_45156# AVSS 0.00125f $ **FLOATING
C14781 a_920_45156# AVSS 0.00125f $ **FLOATING
C14782 a_n232_45156# AVSS 0.366f $ **FLOATING
C14783 XA8.XA1.XA5.MN2.D AVSS 2.5f
C14784 XA7.XA1.XA5.MN2.D AVSS 2.49f
C14785 XA6.XA1.XA5.MN2.D AVSS 2.49f
C14786 XA5.XA1.XA5.MN2.D AVSS 2.49f
C14787 XA4.XA1.XA5.MN2.D AVSS 2.48f
C14788 XA3.XA1.XA5.MN2.D AVSS 2.47f
C14789 XA2.XA1.XA5.MN2.D AVSS 2.47f
C14790 XA1.XA1.XA5.MN2.D AVSS 2.46f
C14791 XA0.XA1.XA5.MN2.D AVSS 2.48f
C14792 a_23600_45508# AVSS 0.363f $ **FLOATING
C14793 a_22448_45508# AVSS 0.00152f $ **FLOATING
C14794 a_21080_45508# AVSS 0.00152f $ **FLOATING
C14795 a_19928_45508# AVSS 0.405f $ **FLOATING
C14796 a_18560_45508# AVSS 0.405f $ **FLOATING
C14797 a_17408_45508# AVSS 0.00125f $ **FLOATING
C14798 a_16040_45508# AVSS 0.00125f $ **FLOATING
C14799 a_14888_45508# AVSS 0.405f $ **FLOATING
C14800 a_13520_45508# AVSS 0.405f $ **FLOATING
C14801 a_12368_45508# AVSS 0.00125f $ **FLOATING
C14802 a_11000_45508# AVSS 0.00125f $ **FLOATING
C14803 a_9848_45508# AVSS 0.405f $ **FLOATING
C14804 a_8480_45508# AVSS 0.404f $ **FLOATING
C14805 a_7328_45508# AVSS 0.00125f $ **FLOATING
C14806 a_5960_45508# AVSS 0.00125f $ **FLOATING
C14807 a_4808_45508# AVSS 0.404f $ **FLOATING
C14808 a_3440_45508# AVSS 0.403f $ **FLOATING
C14809 a_2288_45508# AVSS 0.00125f $ **FLOATING
C14810 a_920_45508# AVSS 0.00125f $ **FLOATING
C14811 a_n232_45508# AVSS 0.405f $ **FLOATING
C14812 a_23600_45860# AVSS 0.404f $ **FLOATING
C14813 a_22448_45860# AVSS 0.00152f $ **FLOATING
C14814 a_21080_45860# AVSS 0.00129f $ **FLOATING
C14815 a_19928_45860# AVSS 0.366f $ **FLOATING
C14816 a_18560_45860# AVSS 0.366f $ **FLOATING
C14817 a_17408_45860# AVSS 0.00125f $ **FLOATING
C14818 a_16040_45860# AVSS 0.00125f $ **FLOATING
C14819 a_14888_45860# AVSS 0.366f $ **FLOATING
C14820 a_13520_45860# AVSS 0.366f $ **FLOATING
C14821 a_12368_45860# AVSS 0.00125f $ **FLOATING
C14822 a_11000_45860# AVSS 0.00125f $ **FLOATING
C14823 a_9848_45860# AVSS 0.366f $ **FLOATING
C14824 a_8480_45860# AVSS 0.366f $ **FLOATING
C14825 a_7328_45860# AVSS 0.00125f $ **FLOATING
C14826 a_5960_45860# AVSS 0.00125f $ **FLOATING
C14827 a_4808_45860# AVSS 0.366f $ **FLOATING
C14828 a_3440_45860# AVSS 0.366f $ **FLOATING
C14829 a_2288_45860# AVSS 0.00125f $ **FLOATING
C14830 a_920_45860# AVSS 0.00125f $ **FLOATING
C14831 a_n232_45860# AVSS 0.366f $ **FLOATING
C14832 a_23600_46212# AVSS 0.368f $ **FLOATING
C14833 a_22448_46212# AVSS 0.00152f $ **FLOATING
C14834 a_21080_46212# AVSS 0.00152f $ **FLOATING
C14835 a_19928_46212# AVSS 0.415f $ **FLOATING
C14836 a_18560_46212# AVSS 0.415f $ **FLOATING
C14837 a_17408_46212# AVSS 0.00125f $ **FLOATING
C14838 a_16040_46212# AVSS 0.00125f $ **FLOATING
C14839 a_14888_46212# AVSS 0.415f $ **FLOATING
C14840 a_13520_46212# AVSS 0.415f $ **FLOATING
C14841 a_12368_46212# AVSS 0.00125f $ **FLOATING
C14842 a_11000_46212# AVSS 0.00125f $ **FLOATING
C14843 a_9848_46212# AVSS 0.415f $ **FLOATING
C14844 a_8480_46212# AVSS 0.415f $ **FLOATING
C14845 a_7328_46212# AVSS 0.00125f $ **FLOATING
C14846 a_5960_46212# AVSS 0.00125f $ **FLOATING
C14847 a_4808_46212# AVSS 0.415f $ **FLOATING
C14848 a_3440_46212# AVSS 0.415f $ **FLOATING
C14849 a_2288_46212# AVSS 0.00125f $ **FLOATING
C14850 a_920_46212# AVSS 0.00125f $ **FLOATING
C14851 a_n232_46212# AVSS 0.416f $ **FLOATING
C14852 XA20.XA2a.MN0.D AVSS 17.9f
C14853 a_23600_46564# AVSS 0.404f $ **FLOATING
C14854 a_22448_46564# AVSS 0.00152f $ **FLOATING
C14855 a_21080_46564# AVSS 0.00152f $ **FLOATING
C14856 a_19928_46564# AVSS 0.366f $ **FLOATING
C14857 a_18560_46564# AVSS 0.366f $ **FLOATING
C14858 a_17408_46564# AVSS 0.00125f $ **FLOATING
C14859 a_16040_46564# AVSS 0.00125f $ **FLOATING
C14860 a_14888_46564# AVSS 0.366f $ **FLOATING
C14861 a_13520_46564# AVSS 0.366f $ **FLOATING
C14862 a_12368_46564# AVSS 0.00125f $ **FLOATING
C14863 a_11000_46564# AVSS 0.00125f $ **FLOATING
C14864 a_9848_46564# AVSS 0.366f $ **FLOATING
C14865 a_8480_46564# AVSS 0.366f $ **FLOATING
C14866 a_7328_46564# AVSS 0.00125f $ **FLOATING
C14867 a_5960_46564# AVSS 0.00125f $ **FLOATING
C14868 a_4808_46564# AVSS 0.366f $ **FLOATING
C14869 a_3440_46564# AVSS 0.366f $ **FLOATING
C14870 a_2288_46564# AVSS 0.00125f $ **FLOATING
C14871 a_920_46564# AVSS 0.00125f $ **FLOATING
C14872 a_n232_46564# AVSS 0.366f $ **FLOATING
C14873 XA8.XA3.MN0.G AVSS 3.68f
C14874 XA7.XA3.MN0.G AVSS 3.66f
C14875 XA6.XA3.MN0.G AVSS 3.66f
C14876 XA5.XA3.MN0.G AVSS 3.66f
C14877 XA4.XA3.MN0.G AVSS 3.66f
C14878 XA3.XA3.MN0.G AVSS 11f
C14879 XA2.XA3.MN0.G AVSS 11.1f
C14880 XA1.XA3.MN0.G AVSS 10.4f
C14881 D<8> AVSS 19.5f
C14882 a_23600_46916# AVSS 0.368f $ **FLOATING
C14883 a_22448_46916# AVSS 0.00152f $ **FLOATING
C14884 a_21080_46916# AVSS 0.00159f $ **FLOATING
C14885 a_19928_46916# AVSS 0.406f $ **FLOATING
C14886 a_18560_46916# AVSS 0.406f $ **FLOATING
C14887 a_17408_46916# AVSS 0.00131f $ **FLOATING
C14888 a_16040_46916# AVSS 0.00131f $ **FLOATING
C14889 a_14888_46916# AVSS 0.406f $ **FLOATING
C14890 a_13520_46916# AVSS 0.406f $ **FLOATING
C14891 a_12368_46916# AVSS 0.00131f $ **FLOATING
C14892 a_11000_46916# AVSS 0.00131f $ **FLOATING
C14893 a_9848_46916# AVSS 0.406f $ **FLOATING
C14894 a_8480_46916# AVSS 0.406f $ **FLOATING
C14895 a_7328_46916# AVSS 0.00131f $ **FLOATING
C14896 a_5960_46916# AVSS 0.00131f $ **FLOATING
C14897 a_4808_46916# AVSS 0.406f $ **FLOATING
C14898 a_3440_46916# AVSS 0.406f $ **FLOATING
C14899 a_2288_46916# AVSS 0.00131f $ **FLOATING
C14900 a_920_46916# AVSS 0.00131f $ **FLOATING
C14901 a_n232_46916# AVSS 0.406f $ **FLOATING
C14902 a_23600_47268# AVSS 0.404f $ **FLOATING
C14903 a_22448_47268# AVSS 0.00152f $ **FLOATING
C14904 a_21080_47268# AVSS 0.00129f $ **FLOATING
C14905 a_19928_47268# AVSS 0.366f $ **FLOATING
C14906 a_18560_47268# AVSS 0.366f $ **FLOATING
C14907 a_17408_47268# AVSS 0.00125f $ **FLOATING
C14908 a_16040_47268# AVSS 0.00125f $ **FLOATING
C14909 a_14888_47268# AVSS 0.366f $ **FLOATING
C14910 a_13520_47268# AVSS 0.366f $ **FLOATING
C14911 a_12368_47268# AVSS 0.00125f $ **FLOATING
C14912 a_11000_47268# AVSS 0.00125f $ **FLOATING
C14913 a_9848_47268# AVSS 0.366f $ **FLOATING
C14914 a_8480_47268# AVSS 0.366f $ **FLOATING
C14915 a_7328_47268# AVSS 0.00125f $ **FLOATING
C14916 a_5960_47268# AVSS 0.00125f $ **FLOATING
C14917 a_4808_47268# AVSS 0.366f $ **FLOATING
C14918 a_3440_47268# AVSS 0.366f $ **FLOATING
C14919 a_2288_47268# AVSS 0.00125f $ **FLOATING
C14920 a_920_47268# AVSS 0.00125f $ **FLOATING
C14921 a_n232_47268# AVSS 0.366f $ **FLOATING
C14922 a_23600_47620# AVSS 0.368f $ **FLOATING
C14923 a_22448_47620# AVSS 0.00152f $ **FLOATING
C14924 a_21080_47620# AVSS 0.00152f $ **FLOATING
C14925 a_19928_47620# AVSS 0.414f $ **FLOATING
C14926 a_18560_47620# AVSS 0.414f $ **FLOATING
C14927 a_17408_47620# AVSS 0.00125f $ **FLOATING
C14928 a_16040_47620# AVSS 0.00125f $ **FLOATING
C14929 a_14888_47620# AVSS 0.414f $ **FLOATING
C14930 a_13520_47620# AVSS 0.414f $ **FLOATING
C14931 a_12368_47620# AVSS 0.00125f $ **FLOATING
C14932 a_11000_47620# AVSS 0.00125f $ **FLOATING
C14933 a_9848_47620# AVSS 0.414f $ **FLOATING
C14934 a_8480_47620# AVSS 0.414f $ **FLOATING
C14935 a_7328_47620# AVSS 0.00125f $ **FLOATING
C14936 a_5960_47620# AVSS 0.00125f $ **FLOATING
C14937 a_4808_47620# AVSS 0.414f $ **FLOATING
C14938 a_3440_47620# AVSS 0.414f $ **FLOATING
C14939 a_2288_47620# AVSS 0.00125f $ **FLOATING
C14940 a_920_47620# AVSS 0.00125f $ **FLOATING
C14941 a_n232_47620# AVSS 0.414f $ **FLOATING
C14942 XA20.XA3a.MN0.D AVSS 22.7f
C14943 a_23600_47972# AVSS 0.404f $ **FLOATING
C14944 a_22448_47972# AVSS 0.00152f $ **FLOATING
C14945 a_21080_47972# AVSS 0.00152f $ **FLOATING
C14946 a_19928_47972# AVSS 0.366f $ **FLOATING
C14947 a_18560_47972# AVSS 0.366f $ **FLOATING
C14948 a_17408_47972# AVSS 0.00125f $ **FLOATING
C14949 a_16040_47972# AVSS 0.00125f $ **FLOATING
C14950 a_14888_47972# AVSS 0.366f $ **FLOATING
C14951 a_13520_47972# AVSS 0.366f $ **FLOATING
C14952 a_12368_47972# AVSS 0.00125f $ **FLOATING
C14953 a_11000_47972# AVSS 0.00125f $ **FLOATING
C14954 a_9848_47972# AVSS 0.366f $ **FLOATING
C14955 a_8480_47972# AVSS 0.366f $ **FLOATING
C14956 a_7328_47972# AVSS 0.00125f $ **FLOATING
C14957 a_5960_47972# AVSS 0.00125f $ **FLOATING
C14958 a_4808_47972# AVSS 0.366f $ **FLOATING
C14959 a_3440_47972# AVSS 0.366f $ **FLOATING
C14960 a_2288_47972# AVSS 0.00125f $ **FLOATING
C14961 a_920_47972# AVSS 0.00125f $ **FLOATING
C14962 a_n232_47972# AVSS 0.366f $ **FLOATING
C14963 XA8.XA4.MN0.G AVSS 3.84f
C14964 XA7.XA4.MN0.G AVSS 3.82f
C14965 XA6.XA4.MN0.G AVSS 3.82f
C14966 XA5.XA4.MN0.G AVSS 3.82f
C14967 XA4.XA4.MN0.G AVSS 3.82f
C14968 XA3.XA4.MN0.G AVSS 3.81f
C14969 XA2.XA4.MN0.G AVSS 3.82f
C14970 XA1.XA4.MN0.G AVSS 3.81f
C14971 XA0.XA4.MN0.G AVSS 3.96f
C14972 a_23600_48324# AVSS 0.362f $ **FLOATING
C14973 a_22448_48324# AVSS 0.00152f $ **FLOATING
C14974 a_21080_48324# AVSS 0.00152f $ **FLOATING
C14975 a_19928_48324# AVSS 0.405f $ **FLOATING
C14976 a_18560_48324# AVSS 0.405f $ **FLOATING
C14977 a_17408_48324# AVSS 0.00125f $ **FLOATING
C14978 a_16040_48324# AVSS 0.00125f $ **FLOATING
C14979 a_14888_48324# AVSS 0.405f $ **FLOATING
C14980 a_13520_48324# AVSS 0.405f $ **FLOATING
C14981 a_12368_48324# AVSS 0.00125f $ **FLOATING
C14982 a_11000_48324# AVSS 0.00125f $ **FLOATING
C14983 a_9848_48324# AVSS 0.405f $ **FLOATING
C14984 a_8480_48324# AVSS 0.405f $ **FLOATING
C14985 a_7328_48324# AVSS 0.00125f $ **FLOATING
C14986 a_5960_48324# AVSS 0.00125f $ **FLOATING
C14987 a_4808_48324# AVSS 0.405f $ **FLOATING
C14988 a_3440_48324# AVSS 0.405f $ **FLOATING
C14989 a_2288_48324# AVSS 0.00125f $ **FLOATING
C14990 a_920_48324# AVSS 0.00125f $ **FLOATING
C14991 a_n232_48324# AVSS 0.405f $ **FLOATING
C14992 a_23600_48676# AVSS 0.358f $ **FLOATING
C14993 a_22448_48676# AVSS 0.00152f $ **FLOATING
C14994 a_21080_48676# AVSS 0.00129f $ **FLOATING
C14995 a_19928_48676# AVSS 0.366f $ **FLOATING
C14996 a_18560_48676# AVSS 0.366f $ **FLOATING
C14997 a_17408_48676# AVSS 0.00129f $ **FLOATING
C14998 a_16040_48676# AVSS 0.00129f $ **FLOATING
C14999 a_14888_48676# AVSS 0.366f $ **FLOATING
C15000 a_13520_48676# AVSS 0.366f $ **FLOATING
C15001 a_12368_48676# AVSS 0.00129f $ **FLOATING
C15002 a_11000_48676# AVSS 0.00129f $ **FLOATING
C15003 a_9848_48676# AVSS 0.366f $ **FLOATING
C15004 a_8480_48676# AVSS 0.366f $ **FLOATING
C15005 a_7328_48676# AVSS 0.00129f $ **FLOATING
C15006 a_5960_48676# AVSS 0.00129f $ **FLOATING
C15007 a_4808_48676# AVSS 0.366f $ **FLOATING
C15008 a_3440_48676# AVSS 0.366f $ **FLOATING
C15009 a_2288_48676# AVSS 0.00129f $ **FLOATING
C15010 a_920_48676# AVSS 0.00129f $ **FLOATING
C15011 a_n232_48676# AVSS 0.366f $ **FLOATING
C15012 a_23600_49028# AVSS 0.357f $ **FLOATING
C15013 a_22448_49028# AVSS 0.00152f $ **FLOATING
C15014 a_21080_49028# AVSS 0.00152f $ **FLOATING
C15015 a_19928_49028# AVSS 0.416f $ **FLOATING
C15016 a_18560_49028# AVSS 0.416f $ **FLOATING
C15017 a_17408_49028# AVSS 0.00152f $ **FLOATING
C15018 a_16040_49028# AVSS 0.00152f $ **FLOATING
C15019 a_14888_49028# AVSS 0.416f $ **FLOATING
C15020 a_13520_49028# AVSS 0.416f $ **FLOATING
C15021 a_12368_49028# AVSS 0.00152f $ **FLOATING
C15022 a_11000_49028# AVSS 0.00152f $ **FLOATING
C15023 a_9848_49028# AVSS 0.416f $ **FLOATING
C15024 a_8480_49028# AVSS 0.416f $ **FLOATING
C15025 a_7328_49028# AVSS 0.00152f $ **FLOATING
C15026 a_5960_49028# AVSS 0.00152f $ **FLOATING
C15027 a_4808_49028# AVSS 0.416f $ **FLOATING
C15028 a_3440_49028# AVSS 0.416f $ **FLOATING
C15029 a_2288_49028# AVSS 0.00152f $ **FLOATING
C15030 a_920_49028# AVSS 0.00152f $ **FLOATING
C15031 a_n232_49028# AVSS 0.416f $ **FLOATING
C15032 a_23600_49380# AVSS 0.357f $ **FLOATING
C15033 a_22448_49380# AVSS 0.00148f $ **FLOATING
C15034 a_21080_49380# AVSS 0.00152f $ **FLOATING
C15035 a_19928_49380# AVSS 0.366f $ **FLOATING
C15036 a_18560_49380# AVSS 0.366f $ **FLOATING
C15037 a_17408_49380# AVSS 0.00152f $ **FLOATING
C15038 a_16040_49380# AVSS 0.00152f $ **FLOATING
C15039 a_14888_49380# AVSS 0.366f $ **FLOATING
C15040 a_13520_49380# AVSS 0.366f $ **FLOATING
C15041 a_12368_49380# AVSS 0.00152f $ **FLOATING
C15042 a_11000_49380# AVSS 0.00152f $ **FLOATING
C15043 a_9848_49380# AVSS 0.366f $ **FLOATING
C15044 a_8480_49380# AVSS 0.366f $ **FLOATING
C15045 a_7328_49380# AVSS 0.00152f $ **FLOATING
C15046 a_5960_49380# AVSS 0.00152f $ **FLOATING
C15047 a_4808_49380# AVSS 0.366f $ **FLOATING
C15048 a_3440_49380# AVSS 0.366f $ **FLOATING
C15049 a_2288_49380# AVSS 0.00152f $ **FLOATING
C15050 a_920_49380# AVSS 0.00152f $ **FLOATING
C15051 a_n232_49380# AVSS 0.366f $ **FLOATING
C15052 XA8.XA4.MN0.D AVSS 3.72f
C15053 XA7.XA4.MN0.D AVSS 3.72f
C15054 XA6.XA4.MN0.D AVSS 3.72f
C15055 XA5.XA4.MN0.D AVSS 3.72f
C15056 XA4.XA4.MN0.D AVSS 3.72f
C15057 XA3.XA4.MN0.D AVSS 6.94f
C15058 XA2.XA4.MN0.D AVSS 7.16f
C15059 XA1.XA4.MN0.D AVSS 12.6f
C15060 VREF AVSS 27.8f
C15061 XA0.XA4.MN0.D AVSS 17.3f
C15062 a_23600_49732# AVSS 0.358f $ **FLOATING
C15063 a_22448_49732# AVSS 0.00148f $ **FLOATING
C15064 a_21080_49732# AVSS 0.00159f $ **FLOATING
C15065 a_19928_49732# AVSS 0.406f $ **FLOATING
C15066 a_18560_49732# AVSS 0.406f $ **FLOATING
C15067 a_17408_49732# AVSS 0.00159f $ **FLOATING
C15068 a_16040_49732# AVSS 0.00159f $ **FLOATING
C15069 a_14888_49732# AVSS 0.406f $ **FLOATING
C15070 a_13520_49732# AVSS 0.406f $ **FLOATING
C15071 a_12368_49732# AVSS 0.00159f $ **FLOATING
C15072 a_11000_49732# AVSS 0.00159f $ **FLOATING
C15073 a_9848_49732# AVSS 0.406f $ **FLOATING
C15074 a_8480_49732# AVSS 0.406f $ **FLOATING
C15075 a_7328_49732# AVSS 0.00159f $ **FLOATING
C15076 a_5960_49732# AVSS 0.00159f $ **FLOATING
C15077 a_4808_49732# AVSS 0.406f $ **FLOATING
C15078 a_3440_49732# AVSS 0.406f $ **FLOATING
C15079 a_2288_49732# AVSS 0.00159f $ **FLOATING
C15080 a_920_49732# AVSS 0.00159f $ **FLOATING
C15081 a_n232_49732# AVSS 0.406f $ **FLOATING
C15082 XA20.XA3.MN0.D AVSS 2.31f
C15083 a_23600_50084# AVSS 0.359f $ **FLOATING
C15084 a_22448_50084# AVSS 0.00148f $ **FLOATING
C15085 a_21080_50084# AVSS 0.00152f $ **FLOATING
C15086 a_19928_50084# AVSS 0.366f $ **FLOATING
C15087 a_18560_50084# AVSS 0.363f $ **FLOATING
C15088 a_17408_50084# AVSS 0.00143f $ **FLOATING
C15089 a_16040_50084# AVSS 0.00143f $ **FLOATING
C15090 a_14888_50084# AVSS 0.363f $ **FLOATING
C15091 a_13520_50084# AVSS 0.363f $ **FLOATING
C15092 a_12368_50084# AVSS 0.00143f $ **FLOATING
C15093 a_11000_50084# AVSS 0.00143f $ **FLOATING
C15094 a_9848_50084# AVSS 0.363f $ **FLOATING
C15095 a_8480_50084# AVSS 0.363f $ **FLOATING
C15096 a_7328_50084# AVSS 0.00143f $ **FLOATING
C15097 a_5960_50084# AVSS 0.00143f $ **FLOATING
C15098 a_4808_50084# AVSS 0.363f $ **FLOATING
C15099 a_3440_50084# AVSS 0.363f $ **FLOATING
C15100 a_2288_50084# AVSS 0.00143f $ **FLOATING
C15101 a_920_50084# AVSS 0.00143f $ **FLOATING
C15102 a_n232_50084# AVSS 0.363f $ **FLOATING
C15103 XA20.XA3.MN1.D AVSS 0.597f
C15104 XA20.XA3.MN6.D AVSS 3.02f
C15105 XA20.XA3a.MN0.G AVSS 2.98f
C15106 XA8.XA6.MP0.D AVSS 0.00592f
C15107 XA8.XA6.MN0.D AVSS 0.218f
C15108 XA8.XA6.MP0.G AVSS 0.964f
C15109 XA7.XA6.MN0.D AVSS 0.201f
C15110 XA7.XA6.MP0.D AVSS 0.00592f
C15111 XA7.XA6.MP0.G AVSS 8.77f
C15112 XA6.XA6.MP0.D AVSS 0.00592f
C15113 XA6.XA6.MN0.D AVSS 0.201f
C15114 XA6.XA6.MP0.G AVSS 6.39f
C15115 XA5.XA6.MN0.D AVSS 0.201f
C15116 XA5.XA6.MP0.D AVSS 0.00592f
C15117 XA5.XA6.MP0.G AVSS 5.21f
C15118 XA4.XA6.MP0.D AVSS 0.00592f
C15119 XA4.XA6.MN0.D AVSS 0.201f
C15120 XA4.XA6.MP0.G AVSS 6.53f
C15121 XA3.XA6.MN0.D AVSS 0.201f
C15122 XA3.XA6.MP0.D AVSS 0.00592f
C15123 XA3.XA6.MP0.G AVSS 4.62f
C15124 XA2.XA6.MP0.D AVSS 0.00592f
C15125 XA2.XA6.MN0.D AVSS 0.201f
C15126 XA2.XA6.MP0.G AVSS 4.95f
C15127 XA1.XA6.MN0.D AVSS 0.201f
C15128 XA1.XA6.MP0.D AVSS 0.00592f
C15129 XA1.XA6.MP0.G AVSS 10.5f
C15130 XA0.XA6.MP0.D AVSS 0.00592f
C15131 XA0.XA6.MN0.D AVSS 0.201f
C15132 XA0.XA6.MP0.G AVSS 15.1f
C15133 a_23600_50436# AVSS 0.381f $ **FLOATING
C15134 a_22448_50436# AVSS 0.00152f $ **FLOATING
C15135 a_21080_50436# AVSS 0.00152f $ **FLOATING
C15136 a_19928_50436# AVSS 0.416f $ **FLOATING
C15137 a_18560_50436# AVSS 0.415f $ **FLOATING
C15138 a_17408_50436# AVSS 0.00152f $ **FLOATING
C15139 a_16040_50436# AVSS 0.00152f $ **FLOATING
C15140 a_14888_50436# AVSS 0.415f $ **FLOATING
C15141 a_13520_50436# AVSS 0.415f $ **FLOATING
C15142 a_12368_50436# AVSS 0.00152f $ **FLOATING
C15143 a_11000_50436# AVSS 0.00152f $ **FLOATING
C15144 a_9848_50436# AVSS 0.415f $ **FLOATING
C15145 a_8480_50436# AVSS 0.415f $ **FLOATING
C15146 a_7328_50436# AVSS 0.00152f $ **FLOATING
C15147 a_5960_50436# AVSS 0.00152f $ **FLOATING
C15148 a_4808_50436# AVSS 0.415f $ **FLOATING
C15149 a_3440_50436# AVSS 0.415f $ **FLOATING
C15150 a_2288_50436# AVSS 0.00152f $ **FLOATING
C15151 a_920_50436# AVSS 0.00152f $ **FLOATING
C15152 a_n232_50436# AVSS 0.416f $ **FLOATING
C15153 a_23600_50788# AVSS 0.361f $ **FLOATING
C15154 a_22448_50788# AVSS 0.00152f $ **FLOATING
C15155 a_21080_50788# AVSS 0.00152f $ **FLOATING
C15156 a_19928_50788# AVSS 0.361f $ **FLOATING
C15157 a_18560_50788# AVSS 0.363f $ **FLOATING
C15158 a_17408_50788# AVSS 0.00152f $ **FLOATING
C15159 a_16040_50788# AVSS 0.00152f $ **FLOATING
C15160 a_14888_50788# AVSS 0.363f $ **FLOATING
C15161 a_13520_50788# AVSS 0.363f $ **FLOATING
C15162 a_12368_50788# AVSS 0.00152f $ **FLOATING
C15163 a_11000_50788# AVSS 0.00152f $ **FLOATING
C15164 a_9848_50788# AVSS 0.363f $ **FLOATING
C15165 a_8480_50788# AVSS 0.363f $ **FLOATING
C15166 a_7328_50788# AVSS 0.00152f $ **FLOATING
C15167 a_5960_50788# AVSS 0.00152f $ **FLOATING
C15168 a_4808_50788# AVSS 0.363f $ **FLOATING
C15169 a_3440_50788# AVSS 0.363f $ **FLOATING
C15170 a_2288_50788# AVSS 0.00152f $ **FLOATING
C15171 a_920_50788# AVSS 0.00152f $ **FLOATING
C15172 a_n232_50788# AVSS 0.363f $ **FLOATING
C15173 XA8.XA6.MP2.D AVSS 0.00592f
C15174 XA8.XA6.MN2.D AVSS 0.141f
C15175 D<0> AVSS 1.24f
C15176 XA7.XA6.MN2.D AVSS 0.15f
C15177 XA7.XA6.MP2.D AVSS 0.00592f
C15178 D<1> AVSS 11.9f
C15179 XA6.XA6.MP2.D AVSS 0.00592f
C15180 XA6.XA6.MN2.D AVSS 0.15f
C15181 D<2> AVSS 9.38f
C15182 XA5.XA6.MN2.D AVSS 0.15f
C15183 XA5.XA6.MP2.D AVSS 0.00592f
C15184 D<3> AVSS 8.3f
C15185 XA4.XA6.MP2.D AVSS 0.00592f
C15186 XA4.XA6.MN2.D AVSS 0.15f
C15187 D<4> AVSS 8.94f
C15188 XA3.XA6.MN2.D AVSS 0.15f
C15189 XA3.XA6.MP2.D AVSS 0.00592f
C15190 D<5> AVSS 8.41f
C15191 XA2.XA6.MP2.D AVSS 0.00592f
C15192 XA2.XA6.MN2.D AVSS 0.15f
C15193 D<6> AVSS 9.41f
C15194 XA1.XA6.MN2.D AVSS 0.15f
C15195 XA1.XA6.MP2.D AVSS 0.00592f
C15196 D<7> AVSS 8.44f
C15197 XA0.XA6.MP2.D AVSS 0.00592f
C15198 XA0.XA6.MN2.D AVSS 0.15f
C15199 XA0.XA6.MP2.G AVSS 14.9f
C15200 a_23600_51140# AVSS 0.358f $ **FLOATING
C15201 a_22448_51140# AVSS 0.00152f $ **FLOATING
C15202 a_21080_51140# AVSS 0.00159f $ **FLOATING
C15203 a_19928_51140# AVSS 0.382f $ **FLOATING
C15204 a_18560_51140# AVSS 0.383f $ **FLOATING
C15205 a_17408_51140# AVSS 0.00159f $ **FLOATING
C15206 a_16040_51140# AVSS 0.00159f $ **FLOATING
C15207 a_14888_51140# AVSS 0.383f $ **FLOATING
C15208 a_13520_51140# AVSS 0.383f $ **FLOATING
C15209 a_12368_51140# AVSS 0.00159f $ **FLOATING
C15210 a_11000_51140# AVSS 0.00159f $ **FLOATING
C15211 a_9848_51140# AVSS 0.383f $ **FLOATING
C15212 a_8480_51140# AVSS 0.383f $ **FLOATING
C15213 a_7328_51140# AVSS 0.00159f $ **FLOATING
C15214 a_5960_51140# AVSS 0.00159f $ **FLOATING
C15215 a_4808_51140# AVSS 0.383f $ **FLOATING
C15216 a_3440_51140# AVSS 0.383f $ **FLOATING
C15217 a_2288_51140# AVSS 0.00159f $ **FLOATING
C15218 a_920_51140# AVSS 0.00159f $ **FLOATING
C15219 a_n232_51140# AVSS 0.383f $ **FLOATING
C15220 XA8.XA7.MP0.G AVSS 1.85f
C15221 XA8.XA1.XA5.MN2.G AVSS 4.7f
C15222 XA7.XA1.XA5.MN2.G AVSS 4.58f
C15223 XA6.XA1.XA5.MN2.G AVSS 4.65f
C15224 XA5.XA1.XA5.MN2.G AVSS 4.59f
C15225 XA4.XA1.XA5.MN2.G AVSS 4.67f
C15226 XA3.XA1.XA5.MN2.G AVSS 4.64f
C15227 XA2.XA1.XA5.MN2.G AVSS 4.63f
C15228 XA0.XA7.MP0.G AVSS 4.64f
C15229 a_23600_51492# AVSS 0.357f $ **FLOATING
C15230 a_22448_51492# AVSS 0.00152f $ **FLOATING
C15231 a_21080_51492# AVSS 0.00152f $ **FLOATING
C15232 a_19928_51492# AVSS 0.387f $ **FLOATING
C15233 a_18560_51492# AVSS 0.387f $ **FLOATING
C15234 a_17408_51492# AVSS 0.00152f $ **FLOATING
C15235 a_16040_51492# AVSS 0.00152f $ **FLOATING
C15236 a_14888_51492# AVSS 0.387f $ **FLOATING
C15237 a_13520_51492# AVSS 0.387f $ **FLOATING
C15238 a_12368_51492# AVSS 0.00152f $ **FLOATING
C15239 a_11000_51492# AVSS 0.00152f $ **FLOATING
C15240 a_9848_51492# AVSS 0.387f $ **FLOATING
C15241 a_8480_51492# AVSS 0.387f $ **FLOATING
C15242 a_7328_51492# AVSS 0.00152f $ **FLOATING
C15243 a_5960_51492# AVSS 0.00152f $ **FLOATING
C15244 a_4808_51492# AVSS 0.387f $ **FLOATING
C15245 a_3440_51492# AVSS 0.387f $ **FLOATING
C15246 a_2288_51492# AVSS 0.00152f $ **FLOATING
C15247 a_920_51492# AVSS 0.00152f $ **FLOATING
C15248 a_n232_51492# AVSS 0.388f $ **FLOATING
C15249 XA7.XA8.MP0.D AVSS 0.223f
C15250 XA6.XA8.MP0.D AVSS 0.223f
C15251 XA5.XA8.MP0.D AVSS 0.223f
C15252 XA4.XA8.MP0.D AVSS 0.223f
C15253 XA3.XA8.MP0.D AVSS 0.223f
C15254 XA2.XA8.MP0.D AVSS 0.223f
C15255 XA1.XA8.MP0.D AVSS 0.223f
C15256 XA0.XA8.MP0.D AVSS 0.223f
C15257 a_23600_51844# AVSS 0.357f $ **FLOATING
C15258 a_22448_51844# AVSS 0.00152f $ **FLOATING
C15259 a_21080_51844# AVSS 0.00152f $ **FLOATING
C15260 a_19928_51844# AVSS 0.384f $ **FLOATING
C15261 a_18560_51844# AVSS 0.386f $ **FLOATING
C15262 a_17408_51844# AVSS 0.00152f $ **FLOATING
C15263 a_16040_51844# AVSS 0.00152f $ **FLOATING
C15264 a_14888_51844# AVSS 0.386f $ **FLOATING
C15265 a_13520_51844# AVSS 0.386f $ **FLOATING
C15266 a_12368_51844# AVSS 0.00152f $ **FLOATING
C15267 a_11000_51844# AVSS 0.00152f $ **FLOATING
C15268 a_9848_51844# AVSS 0.386f $ **FLOATING
C15269 a_8480_51844# AVSS 0.386f $ **FLOATING
C15270 a_7328_51844# AVSS 0.00152f $ **FLOATING
C15271 a_5960_51844# AVSS 0.00152f $ **FLOATING
C15272 a_4808_51844# AVSS 0.386f $ **FLOATING
C15273 a_3440_51844# AVSS 0.386f $ **FLOATING
C15274 a_2288_51844# AVSS 0.00152f $ **FLOATING
C15275 a_920_51844# AVSS 0.00152f $ **FLOATING
C15276 a_n232_51844# AVSS 0.386f $ **FLOATING
C15277 XA8.XA7.MP0.D AVSS 1.52f
C15278 XA7.XA7.MP0.D AVSS 1.53f
C15279 XA6.XA7.MP0.D AVSS 1.53f
C15280 XA5.XA7.MP0.D AVSS 1.53f
C15281 XA4.XA7.MP0.D AVSS 1.53f
C15282 XA3.XA7.MP0.D AVSS 1.53f
C15283 XA2.XA7.MP0.D AVSS 1.53f
C15284 XA1.XA7.MP0.D AVSS 1.53f
C15285 XA0.XA7.MP0.D AVSS 1.53f
C15286 a_23600_52196# AVSS 0.357f $ **FLOATING
C15287 a_22448_52196# AVSS 0.00152f $ **FLOATING
C15288 a_21080_52196# AVSS 0.00152f $ **FLOATING
C15289 a_19928_52196# AVSS 0.364f $ **FLOATING
C15290 a_18560_52196# AVSS 0.364f $ **FLOATING
C15291 a_17408_52196# AVSS 0.00152f $ **FLOATING
C15292 a_16040_52196# AVSS 0.00152f $ **FLOATING
C15293 a_14888_52196# AVSS 0.364f $ **FLOATING
C15294 a_13520_52196# AVSS 0.364f $ **FLOATING
C15295 a_12368_52196# AVSS 0.00152f $ **FLOATING
C15296 a_11000_52196# AVSS 0.00152f $ **FLOATING
C15297 a_9848_52196# AVSS 0.364f $ **FLOATING
C15298 a_8480_52196# AVSS 0.364f $ **FLOATING
C15299 a_7328_52196# AVSS 0.00152f $ **FLOATING
C15300 a_5960_52196# AVSS 0.00152f $ **FLOATING
C15301 a_4808_52196# AVSS 0.364f $ **FLOATING
C15302 a_3440_52196# AVSS 0.364f $ **FLOATING
C15303 a_2288_52196# AVSS 0.00152f $ **FLOATING
C15304 a_920_52196# AVSS 0.00152f $ **FLOATING
C15305 a_n232_52196# AVSS 0.365f $ **FLOATING
C15306 SARN AVSS 0.305p
C15307 XA8.XA9.MN0.D AVSS 0.174f
C15308 XA8.XA9.MN1.G AVSS 1.72f
C15309 XA7.XA9.MN0.D AVSS 0.174f
C15310 XA7.XA9.MN1.G AVSS 1.73f
C15311 XA6.XA9.MN0.D AVSS 0.174f
C15312 XA6.XA9.MN1.G AVSS 1.74f
C15313 XA5.XA9.MN0.D AVSS 0.174f
C15314 XA5.XA9.MN1.G AVSS 1.73f
C15315 XA4.XA9.MN0.D AVSS 0.174f
C15316 XA4.XA9.MN1.G AVSS 1.74f
C15317 XA3.XA9.MN0.D AVSS 0.174f
C15318 XA3.XA9.MN1.G AVSS 1.73f
C15319 XA2.XA9.MN0.D AVSS 0.174f
C15320 XA2.XA9.MN1.G AVSS 1.74f
C15321 XA1.XA9.MN0.D AVSS 0.174f
C15322 XA1.XA9.MN1.G AVSS 1.73f
C15323 XA0.XA9.MN0.D AVSS 0.174f
C15324 XA0.XA9.MN1.G AVSS 1.8f
C15325 a_23600_52548# AVSS 0.359f $ **FLOATING
C15326 a_22448_52548# AVSS 0.00152f $ **FLOATING
C15327 a_21080_52548# AVSS 0.00152f $ **FLOATING
C15328 a_19928_52548# AVSS 0.383f $ **FLOATING
C15329 a_18560_52548# AVSS 0.383f $ **FLOATING
C15330 a_17408_52548# AVSS 0.00152f $ **FLOATING
C15331 a_16040_52548# AVSS 0.00152f $ **FLOATING
C15332 a_14888_52548# AVSS 0.383f $ **FLOATING
C15333 a_13520_52548# AVSS 0.383f $ **FLOATING
C15334 a_12368_52548# AVSS 0.00152f $ **FLOATING
C15335 a_11000_52548# AVSS 0.00152f $ **FLOATING
C15336 a_9848_52548# AVSS 0.383f $ **FLOATING
C15337 a_8480_52548# AVSS 0.383f $ **FLOATING
C15338 a_7328_52548# AVSS 0.00152f $ **FLOATING
C15339 a_5960_52548# AVSS 0.00152f $ **FLOATING
C15340 a_4808_52548# AVSS 0.383f $ **FLOATING
C15341 a_3440_52548# AVSS 0.383f $ **FLOATING
C15342 a_2288_52548# AVSS 0.00152f $ **FLOATING
C15343 a_920_52548# AVSS 0.00152f $ **FLOATING
C15344 a_n232_52548# AVSS 0.383f $ **FLOATING
C15345 XA20.XA4.MN0.D AVSS 0.862f
C15346 XA8.XA10.MP0.G AVSS 0.929f
C15347 XA7.XA10.MP0.G AVSS 0.929f
C15348 XA6.XA10.MP0.G AVSS 0.929f
C15349 XA5.XA10.MP0.G AVSS 0.929f
C15350 XA4.XA10.MP0.G AVSS 0.929f
C15351 XA3.XA10.MP0.G AVSS 0.929f
C15352 XA2.XA10.MP0.G AVSS 0.929f
C15353 XA1.XA10.MP0.G AVSS 0.929f
C15354 XA0.XA10.MP0.G AVSS 0.929f
C15355 a_23600_52900# AVSS 0.382f $ **FLOATING
C15356 a_22448_52900# AVSS 0.00152f $ **FLOATING
C15357 a_21080_52900# AVSS 0.00152f $ **FLOATING
C15358 a_19928_52900# AVSS 0.387f $ **FLOATING
C15359 a_18560_52900# AVSS 0.387f $ **FLOATING
C15360 a_17408_52900# AVSS 0.00152f $ **FLOATING
C15361 a_16040_52900# AVSS 0.00152f $ **FLOATING
C15362 a_14888_52900# AVSS 0.387f $ **FLOATING
C15363 a_13520_52900# AVSS 0.387f $ **FLOATING
C15364 a_12368_52900# AVSS 0.00152f $ **FLOATING
C15365 a_11000_52900# AVSS 0.00152f $ **FLOATING
C15366 a_9848_52900# AVSS 0.387f $ **FLOATING
C15367 a_8480_52900# AVSS 0.387f $ **FLOATING
C15368 a_7328_52900# AVSS 0.00152f $ **FLOATING
C15369 a_5960_52900# AVSS 0.00152f $ **FLOATING
C15370 a_4808_52900# AVSS 0.387f $ **FLOATING
C15371 a_3440_52900# AVSS 0.387f $ **FLOATING
C15372 a_2288_52900# AVSS 0.00152f $ **FLOATING
C15373 a_920_52900# AVSS 0.00152f $ **FLOATING
C15374 a_n232_52900# AVSS 0.388f $ **FLOATING
C15375 XA20.XA9.MP0.D AVSS 6.27f
C15376 XA8.XA10.MP0.D AVSS 0.902f
C15377 XA7.XA10.MP0.D AVSS 0.9f
C15378 XA6.XA10.MP0.D AVSS 0.902f
C15379 XA5.XA10.MP0.D AVSS 0.9f
C15380 XA4.XA10.MP0.D AVSS 0.902f
C15381 XA3.XA10.MP0.D AVSS 0.9f
C15382 XA2.XA10.MP0.D AVSS 0.902f
C15383 XA1.XA10.MP0.D AVSS 0.9f
C15384 XA0.XA10.MP0.D AVSS 0.902f
C15385 a_23600_53252# AVSS 0.388f $ **FLOATING
C15386 a_22448_53252# AVSS 0.00159f $ **FLOATING
C15387 a_21080_53252# AVSS 0.00152f $ **FLOATING
C15388 a_19928_53252# AVSS 0.371f $ **FLOATING
C15389 a_18560_53252# AVSS 0.365f $ **FLOATING
C15390 a_17408_53252# AVSS 0.00143f $ **FLOATING
C15391 a_16040_53252# AVSS 0.00152f $ **FLOATING
C15392 a_14888_53252# AVSS 0.371f $ **FLOATING
C15393 a_13520_53252# AVSS 0.365f $ **FLOATING
C15394 a_12368_53252# AVSS 0.00143f $ **FLOATING
C15395 a_11000_53252# AVSS 0.00152f $ **FLOATING
C15396 a_9848_53252# AVSS 0.371f $ **FLOATING
C15397 a_8480_53252# AVSS 0.365f $ **FLOATING
C15398 a_7328_53252# AVSS 0.00143f $ **FLOATING
C15399 a_5960_53252# AVSS 0.00152f $ **FLOATING
C15400 a_4808_53252# AVSS 0.371f $ **FLOATING
C15401 a_3440_53252# AVSS 0.365f $ **FLOATING
C15402 a_2288_53252# AVSS 0.00143f $ **FLOATING
C15403 a_920_53252# AVSS 0.00152f $ **FLOATING
C15404 a_n232_53252# AVSS 0.371f $ **FLOATING
C15405 XA8.XA11.MP0.D AVSS 0.00597f
C15406 XA7.XA11.MP0.D AVSS 0.00597f
C15407 XA6.XA11.MP0.D AVSS 0.00597f
C15408 XA5.XA11.MP0.D AVSS 0.00597f
C15409 XA4.XA11.MP0.D AVSS 0.00597f
C15410 XA3.XA11.MP0.D AVSS 0.00597f
C15411 XA2.XA11.MP0.D AVSS 0.00597f
C15412 XA1.XA11.MP0.D AVSS 0.00597f
C15413 XA0.XA11.MP0.D AVSS 0.00597f
C15414 XA0.XA11.MN1.G AVSS 42.4f
C15415 a_23600_53604# AVSS 0.363f $ **FLOATING
C15416 a_22448_53604# AVSS 0.00152f $ **FLOATING
C15417 a_21080_53604# AVSS 0.00152f $ **FLOATING
C15418 a_19928_53604# AVSS 0.406f $ **FLOATING
C15419 a_18560_53604# AVSS 0.405f $ **FLOATING
C15420 a_17408_53604# AVSS 0.00152f $ **FLOATING
C15421 a_16040_53604# AVSS 0.00152f $ **FLOATING
C15422 a_14888_53604# AVSS 0.406f $ **FLOATING
C15423 a_13520_53604# AVSS 0.405f $ **FLOATING
C15424 a_12368_53604# AVSS 0.00152f $ **FLOATING
C15425 a_11000_53604# AVSS 0.00152f $ **FLOATING
C15426 a_9848_53604# AVSS 0.406f $ **FLOATING
C15427 a_8480_53604# AVSS 0.405f $ **FLOATING
C15428 a_7328_53604# AVSS 0.00152f $ **FLOATING
C15429 a_5960_53604# AVSS 0.00152f $ **FLOATING
C15430 a_4808_53604# AVSS 0.406f $ **FLOATING
C15431 a_3440_53604# AVSS 0.405f $ **FLOATING
C15432 a_2288_53604# AVSS 0.00152f $ **FLOATING
C15433 a_920_53604# AVSS 0.00152f $ **FLOATING
C15434 a_n232_53604# AVSS 0.406f $ **FLOATING
C15435 XA20.XA10.MN0.D AVSS 0.136f
C15436 XA20.XA10.MN1.D AVSS 7.1f
C15437 XA8.XA12.MP0.G AVSS 1.18f
C15438 XA7.XA12.MP0.G AVSS 1.14f
C15439 XA8.XA11.MN1.G AVSS 1.7f
C15440 XA6.XA12.MP0.G AVSS 1.18f
C15441 XA7.XA11.MN1.G AVSS 1.55f
C15442 XA5.XA12.MP0.G AVSS 1.14f
C15443 XA6.XA11.MN1.G AVSS 1.7f
C15444 XA4.XA12.MP0.G AVSS 1.18f
C15445 XA5.XA11.MN1.G AVSS 1.55f
C15446 XA3.XA12.MP0.G AVSS 1.14f
C15447 XA4.XA11.MN1.G AVSS 1.7f
C15448 XA2.XA12.MP0.G AVSS 1.18f
C15449 XA3.XA11.MN1.G AVSS 1.55f
C15450 XA1.XA12.MP0.G AVSS 1.14f
C15451 XA2.XA11.MN1.G AVSS 1.7f
C15452 XA0.XA12.MP0.G AVSS 1.18f
C15453 XA0.XA12.MP0.D AVSS 1.55f
C15454 a_23600_53956# AVSS 0.383f $ **FLOATING
C15455 a_22448_53956# AVSS 0.00152f $ **FLOATING
C15456 a_21080_53956# AVSS 0.00158f $ **FLOATING
C15457 a_19928_53956# AVSS 0.47f $ **FLOATING
C15458 a_18560_53956# AVSS 0.471f $ **FLOATING
C15459 a_17408_53956# AVSS 0.00159f $ **FLOATING
C15460 a_16040_53956# AVSS 0.00158f $ **FLOATING
C15461 a_14888_53956# AVSS 0.47f $ **FLOATING
C15462 a_13520_53956# AVSS 0.471f $ **FLOATING
C15463 a_12368_53956# AVSS 0.00159f $ **FLOATING
C15464 a_11000_53956# AVSS 0.00158f $ **FLOATING
C15465 a_9848_53956# AVSS 0.47f $ **FLOATING
C15466 a_8480_53956# AVSS 0.471f $ **FLOATING
C15467 a_7328_53956# AVSS 0.00159f $ **FLOATING
C15468 a_5960_53956# AVSS 0.00158f $ **FLOATING
C15469 a_4808_53956# AVSS 0.47f $ **FLOATING
C15470 a_3440_53956# AVSS 0.471f $ **FLOATING
C15471 a_2288_53956# AVSS 0.00159f $ **FLOATING
C15472 a_920_53956# AVSS 0.00158f $ **FLOATING
C15473 a_n232_53956# AVSS 0.47f $ **FLOATING
C15474 CK_SAMPLE AVSS 23.5f
C15475 a_23600_54308# AVSS 0.37f $ **FLOATING
C15476 a_22448_54308# AVSS 0.00152f $ **FLOATING
C15477 a_21080_54308# AVSS 0.0894f $ **FLOATING
C15478 a_19928_54308# AVSS 0.539f $ **FLOATING
C15479 a_18560_54308# AVSS 0.538f $ **FLOATING
C15480 a_17408_54308# AVSS 0.0894f $ **FLOATING
C15481 a_16040_54308# AVSS 0.0894f $ **FLOATING
C15482 a_14888_54308# AVSS 0.539f $ **FLOATING
C15483 a_13520_54308# AVSS 0.538f $ **FLOATING
C15484 a_12368_54308# AVSS 0.0894f $ **FLOATING
C15485 a_11000_54308# AVSS 0.0894f $ **FLOATING
C15486 a_9848_54308# AVSS 0.539f $ **FLOATING
C15487 a_8480_54308# AVSS 0.538f $ **FLOATING
C15488 a_7328_54308# AVSS 0.0894f $ **FLOATING
C15489 a_5960_54308# AVSS 0.0894f $ **FLOATING
C15490 a_4808_54308# AVSS 0.539f $ **FLOATING
C15491 a_3440_54308# AVSS 0.538f $ **FLOATING
C15492 a_2288_54308# AVSS 0.0894f $ **FLOATING
C15493 a_920_54308# AVSS 0.0894f $ **FLOATING
C15494 a_n232_54308# AVSS 0.539f $ **FLOATING
C15495 XA20.XA11.MP0.D AVSS 0.00592f
C15496 DONE AVSS 1.18f
C15497 XA20.XA11.MN0.D AVSS 1.24f
C15498 a_23600_54660# AVSS 0.407f $ **FLOATING
C15499 a_22448_54660# AVSS 0.00276f $ **FLOATING
C15500 XA20.XA12.MP0.G AVSS 1.12f
C15501 XA20.XA12.MP0.D AVSS 0.791f
C15502 a_23600_55012# AVSS 0.471f $ **FLOATING
C15503 a_22448_55012# AVSS 0.00282f $ **FLOATING
C15504 a_23600_55364# AVSS 0.541f $ **FLOATING
C15505 a_22448_55364# AVSS 0.0952f $ **FLOATING
C15506 AVDD AVSS 0.691p
.ends

