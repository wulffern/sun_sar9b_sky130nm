magic
tech sky130A
magscale 1 1
timestamp 1712872800
<< checkpaint >>
rect 0 0 1260 5368
<< locali >>
rect 216 2271 300 2305
rect 300 1875 432 1909
rect 300 1875 334 2305
rect 216 3151 300 3185
rect 300 2755 432 2789
rect 300 2755 334 3185
rect 926 1831 1044 1865
rect 828 1699 926 1733
rect 926 1699 960 1865
rect 216 4207 300 4241
rect 300 4075 432 4109
rect 300 4075 334 4241
rect 199 4207 233 4417
rect 240 4613 300 4647
rect 300 4515 432 4549
rect 300 4515 334 4647
rect 236 4647 270 4681
rect 240 4789 300 4823
rect 300 4691 432 4725
rect 300 4691 334 4823
rect 236 4823 270 4857
rect 216 5087 300 5121
rect 300 4867 432 4901
rect 300 4867 334 5121
rect 828 3195 912 3229
rect 912 3591 1044 3625
rect 912 3195 946 3625
rect 990 1655 1098 1689
rect 162 1479 270 1513
rect 162 4911 270 4945
rect 774 5131 882 5165
rect 162 3679 270 3713
rect 378 4251 486 4285
<< m1 >>
rect 216 2711 300 2745
rect 300 1347 432 1381
rect 300 1347 334 2745
rect 1044 4031 1128 4065
rect 828 379 1128 413
rect 1128 379 1162 4065
rect 216 4471 300 4505
rect 300 3899 432 3933
rect 300 3899 334 4505
rect 828 2315 912 2349
rect 912 3767 1044 3801
rect 912 2315 946 3801
<< m3 >>
rect 1095 1963 1129 3383
rect 170 2269 270 2307
rect 527 2282 565 2382
rect 607 2722 645 2822
rect 695 3162 733 3262
rect 1062 1963 1162 2063
rect 774 0 874 5368
rect 378 0 478 5368
rect 774 0 874 5368
rect 378 0 478 5368
<< m2 >>
rect 178 1127 270 1161
rect 178 247 270 281
rect 790 379 882 413
use SUNSAR_SARMRYX1_CV XA1 
transform 1 0 0 0 1 0
box 0 0 1260 1760
use SUNSAR_SWX4_CV XA2 
transform 1 0 0 0 1 1760
box 0 1760 1260 2200
use SUNSAR_SWX4_CV XA3 
transform 1 0 0 0 1 2200
box 0 2200 1260 2640
use SUNSAR_SWX4_CV XA4 
transform 1 0 0 0 1 2640
box 0 2640 1260 3080
use SUNSAR_SWX4_CV XA5 
transform 1 0 0 0 1 3080
box 0 3080 1260 3520
use SUNSAR_SARCEX1_CV XA6 
transform 1 0 0 0 1 3520
box 0 3520 1260 3960
use SUNSAR_IVX1_CV XA7 
transform 1 0 0 0 1 3960
box 0 3960 1260 4136
use SUNSAR_IVX1_CV XA8 
transform 1 0 0 0 1 4136
box 0 4136 1260 4312
use SUNSAR_NDX1_CV XA9 
transform 1 0 0 0 1 4312
box 0 4312 1260 4576
use SUNSAR_IVX1_CV XA10 
transform 1 0 0 0 1 4576
box 0 4576 1260 4752
use SUNSAR_NRX1_CV XA11 
transform 1 0 0 0 1 4752
box 0 4752 1260 5016
use SUNSAR_IVX1_CV XA12 
transform 1 0 0 0 1 5016
box 0 5016 1260 5192
use SUNSAR_TAPCELLB_CV XA13 
transform 1 0 0 0 1 5192
box 0 5192 1260 5368
use SUNSAR_cut_M1M2_2x1 xcut0 
transform 1 0 162 0 1 2711
box 162 2711 254 2745
use SUNSAR_cut_M1M2_2x1 xcut1 
transform 1 0 378 0 1 1347
box 378 1347 470 1381
use SUNSAR_cut_M1M2_2x1 xcut2 
transform 1 0 990 0 1 4031
box 990 4031 1082 4065
use SUNSAR_cut_M1M2_2x1 xcut3 
transform 1 0 774 0 1 379
box 774 379 866 413
use SUNSAR_cut_M1M2_2x1 xcut4 
transform 1 0 162 0 1 4471
box 162 4471 254 4505
use SUNSAR_cut_M1M2_2x1 xcut5 
transform 1 0 378 0 1 3899
box 378 3899 470 3933
use SUNSAR_cut_M1M2_2x1 xcut6 
transform 1 0 774 0 1 2315
box 774 2315 866 2349
use SUNSAR_cut_M1M2_2x1 xcut7 
transform 1 0 990 0 1 3767
box 990 3767 1082 3801
use SUNSAR_cut_M1M4_2x1 xcut8 
transform 1 0 170 0 1 2269
box 170 2269 270 2307
use SUNSAR_cut_M1M4_1x2 xcut9 
transform 1 0 527 0 1 2282
box 527 2282 565 2382
use SUNSAR_cut_M1M4_1x2 xcut10 
transform 1 0 607 0 1 2722
box 607 2722 645 2822
use SUNSAR_cut_M1M4_1x2 xcut11 
transform 1 0 695 0 1 3162
box 695 3162 733 3262
use SUNSAR_cut_M2M3_2x1 xcut12 
transform 1 0 790 0 1 379
box 790 379 882 413
use SUNSAR_cut_M2M3_2x1 xcut13 
transform 1 0 178 0 1 247
box 178 247 270 281
use SUNSAR_cut_M2M3_2x1 xcut14 
transform 1 0 178 0 1 247
box 178 247 270 281
use SUNSAR_cut_M2M3_2x1 xcut15 
transform 1 0 178 0 1 1127
box 178 1127 270 1161
use SUNSAR_cut_M2M3_2x1 xcut16 
transform 1 0 178 0 1 1127
box 178 1127 270 1161
<< labels >>
flabel m2 s 178 1127 270 1161 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew signal bidirectional
flabel locali s 990 1655 1098 1689 0 FreeSans 400 0 0 0 RST_N
port 4 nsew signal bidirectional
flabel m2 s 178 247 270 281 0 FreeSans 400 0 0 0 EN
port 3 nsew signal bidirectional
flabel locali s 162 1479 270 1513 0 FreeSans 400 0 0 0 CMP_ON
port 2 nsew signal bidirectional
flabel m2 s 790 379 882 413 0 FreeSans 400 0 0 0 ENO
port 5 nsew signal bidirectional
flabel m3 s 170 2269 270 2307 0 FreeSans 400 0 0 0 CN1
port 10 nsew signal bidirectional
flabel m3 s 527 2282 565 2382 0 FreeSans 400 0 0 0 CP1
port 8 nsew signal bidirectional
flabel m3 s 607 2722 645 2822 0 FreeSans 400 0 0 0 CP0
port 7 nsew signal bidirectional
flabel m3 s 695 3162 733 3262 0 FreeSans 400 0 0 0 CN0
port 9 nsew signal bidirectional
flabel locali s 162 4911 270 4945 0 FreeSans 400 0 0 0 CEIN
port 11 nsew signal bidirectional
flabel locali s 774 5131 882 5165 0 FreeSans 400 0 0 0 CEO
port 12 nsew signal bidirectional
flabel locali s 162 3679 270 3713 0 FreeSans 400 0 0 0 CKS
port 13 nsew signal bidirectional
flabel locali s 378 4251 486 4285 0 FreeSans 400 0 0 0 DONE
port 6 nsew signal bidirectional
flabel m3 s 1062 1963 1162 2063 0 FreeSans 400 0 0 0 VREF
port 14 nsew signal bidirectional
flabel m3 s 774 0 874 5368 0 FreeSans 400 0 0 0 AVDD
port 15 nsew signal bidirectional
flabel m3 s 378 0 478 5368 0 FreeSans 400 0 0 0 AVSS
port 16 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 5368
<< end >>
